
module read_sync_addrbits8 ( clk_out, rst, rdptr, sync_rdptr, sync_flush_BAR
 );
  input [8:0] rdptr;
  output [8:0] sync_rdptr;
  input clk_out, rst, sync_flush_BAR;
  wire   sync_flush, N4, N5, N6, N7, N8, N9, N10, N11, N13, N14, N15, N16, N17,
         N18, N19, N20, n1, n2;
  wire   [8:0] r0;
  assign sync_flush = sync_flush_BAR;

  DFFARX1 \r0_reg[7]  ( .D(N11), .CLK(clk_out), .RSTB(rst), .Q(r0[7]) );
  DFFARX1 \r0_reg[6]  ( .D(N10), .CLK(clk_out), .RSTB(rst), .Q(r0[6]) );
  DFFARX1 \r0_reg[5]  ( .D(N9), .CLK(clk_out), .RSTB(rst), .Q(r0[5]) );
  DFFARX1 \r0_reg[4]  ( .D(N8), .CLK(clk_out), .RSTB(rst), .Q(r0[4]) );
  DFFARX1 \r0_reg[3]  ( .D(N7), .CLK(clk_out), .RSTB(n2), .Q(r0[3]) );
  DFFARX1 \r0_reg[2]  ( .D(N6), .CLK(clk_out), .RSTB(n2), .Q(r0[2]) );
  DFFARX1 \r0_reg[1]  ( .D(N5), .CLK(clk_out), .RSTB(n2), .Q(r0[1]) );
  DFFARX1 \r0_reg[0]  ( .D(N4), .CLK(clk_out), .RSTB(n2), .Q(r0[0]) );
  DFFARX1 \sync_rdptr_reg[7]  ( .D(N20), .CLK(clk_out), .RSTB(n2), .Q(
        sync_rdptr[7]) );
  DFFARX1 \sync_rdptr_reg[6]  ( .D(N19), .CLK(clk_out), .RSTB(n2), .Q(
        sync_rdptr[6]) );
  DFFARX1 \sync_rdptr_reg[5]  ( .D(N18), .CLK(clk_out), .RSTB(n2), .Q(
        sync_rdptr[5]) );
  DFFARX1 \sync_rdptr_reg[4]  ( .D(N17), .CLK(clk_out), .RSTB(n2), .Q(
        sync_rdptr[4]) );
  DFFARX1 \sync_rdptr_reg[3]  ( .D(N16), .CLK(clk_out), .RSTB(n2), .Q(
        sync_rdptr[3]) );
  DFFARX1 \sync_rdptr_reg[2]  ( .D(N15), .CLK(clk_out), .RSTB(n2), .Q(
        sync_rdptr[2]) );
  DFFARX1 \sync_rdptr_reg[1]  ( .D(N14), .CLK(clk_out), .RSTB(n2), .Q(
        sync_rdptr[1]) );
  DFFARX1 \sync_rdptr_reg[0]  ( .D(N13), .CLK(clk_out), .RSTB(n2), .Q(
        sync_rdptr[0]) );
  AND2X1 U4 ( .IN1(rdptr[5]), .IN2(sync_flush), .Q(N9) );
  AND2X1 U5 ( .IN1(rdptr[4]), .IN2(n1), .Q(N8) );
  AND2X1 U6 ( .IN1(rdptr[3]), .IN2(n1), .Q(N7) );
  AND2X1 U7 ( .IN1(rdptr[2]), .IN2(n1), .Q(N6) );
  AND2X1 U8 ( .IN1(rdptr[1]), .IN2(sync_flush), .Q(N5) );
  AND2X1 U9 ( .IN1(rdptr[0]), .IN2(n1), .Q(N4) );
  AND2X1 U11 ( .IN1(r0[7]), .IN2(n1), .Q(N20) );
  AND2X1 U12 ( .IN1(r0[6]), .IN2(n1), .Q(N19) );
  AND2X1 U13 ( .IN1(r0[5]), .IN2(sync_flush), .Q(N18) );
  AND2X1 U14 ( .IN1(r0[4]), .IN2(n1), .Q(N17) );
  AND2X1 U15 ( .IN1(r0[3]), .IN2(sync_flush), .Q(N16) );
  AND2X1 U16 ( .IN1(r0[2]), .IN2(n1), .Q(N15) );
  AND2X1 U17 ( .IN1(r0[1]), .IN2(sync_flush), .Q(N14) );
  AND2X1 U18 ( .IN1(r0[0]), .IN2(n1), .Q(N13) );
  AND2X1 U20 ( .IN1(rdptr[7]), .IN2(sync_flush), .Q(N11) );
  AND2X1 U21 ( .IN1(rdptr[6]), .IN2(n1), .Q(N10) );
  NBUFFX2 U3 ( .INP(rst), .Z(n2) );
  NBUFFX2 U10 ( .INP(sync_flush), .Z(n1) );
endmodule


module write_sync_addrbits8 ( clk_in, rst, flush, wrptr, sync_wrptr );
  input [8:0] wrptr;
  output [8:0] sync_wrptr;
  input clk_in, rst, flush;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, n1, n2, n3, n4, n5, n6;
  wire   [8:0] w0;

  DFFARX1 \w0_reg[8]  ( .D(N12), .CLK(clk_in), .RSTB(n5), .QN(n3) );
  DFFARX1 \w0_reg[7]  ( .D(N11), .CLK(clk_in), .RSTB(n5), .QN(n2) );
  DFFARX1 \w0_reg[6]  ( .D(N10), .CLK(clk_in), .RSTB(n5), .QN(n1) );
  DFFARX1 \w0_reg[5]  ( .D(N9), .CLK(clk_in), .RSTB(n5), .Q(w0[5]) );
  DFFARX1 \w0_reg[4]  ( .D(N8), .CLK(clk_in), .RSTB(n5), .Q(w0[4]) );
  DFFARX1 \w0_reg[3]  ( .D(N7), .CLK(clk_in), .RSTB(n5), .Q(w0[3]) );
  DFFARX1 \w0_reg[2]  ( .D(N6), .CLK(clk_in), .RSTB(n4), .Q(w0[2]) );
  DFFARX1 \w0_reg[1]  ( .D(N5), .CLK(clk_in), .RSTB(n4), .Q(w0[1]) );
  DFFARX1 \w0_reg[0]  ( .D(N4), .CLK(clk_in), .RSTB(n4), .Q(w0[0]) );
  DFFARX1 \sync_wrptr_reg[8]  ( .D(N21), .CLK(clk_in), .RSTB(n4), .Q(
        sync_wrptr[8]) );
  DFFARX1 \sync_wrptr_reg[7]  ( .D(N20), .CLK(clk_in), .RSTB(n4), .Q(
        sync_wrptr[7]) );
  DFFARX1 \sync_wrptr_reg[6]  ( .D(N19), .CLK(clk_in), .RSTB(n4), .Q(
        sync_wrptr[6]) );
  DFFARX1 \sync_wrptr_reg[5]  ( .D(N18), .CLK(clk_in), .RSTB(n4), .Q(
        sync_wrptr[5]) );
  DFFARX1 \sync_wrptr_reg[4]  ( .D(N17), .CLK(clk_in), .RSTB(n4), .Q(
        sync_wrptr[4]) );
  DFFARX1 \sync_wrptr_reg[3]  ( .D(N16), .CLK(clk_in), .RSTB(n4), .Q(
        sync_wrptr[3]) );
  DFFARX1 \sync_wrptr_reg[2]  ( .D(N15), .CLK(clk_in), .RSTB(n4), .Q(
        sync_wrptr[2]) );
  DFFARX1 \sync_wrptr_reg[1]  ( .D(N14), .CLK(clk_in), .RSTB(n4), .Q(
        sync_wrptr[1]) );
  DFFARX1 \sync_wrptr_reg[0]  ( .D(N13), .CLK(clk_in), .RSTB(n4), .Q(
        sync_wrptr[0]) );
  AND2X1 U4 ( .IN1(wrptr[5]), .IN2(n6), .Q(N9) );
  AND2X1 U5 ( .IN1(wrptr[4]), .IN2(n6), .Q(N8) );
  AND2X1 U6 ( .IN1(wrptr[3]), .IN2(n6), .Q(N7) );
  AND2X1 U7 ( .IN1(wrptr[2]), .IN2(n6), .Q(N6) );
  AND2X1 U8 ( .IN1(wrptr[1]), .IN2(n6), .Q(N5) );
  AND2X1 U9 ( .IN1(wrptr[0]), .IN2(n6), .Q(N4) );
  AND2X1 U13 ( .IN1(w0[5]), .IN2(n6), .Q(N18) );
  AND2X1 U14 ( .IN1(w0[4]), .IN2(n6), .Q(N17) );
  AND2X1 U15 ( .IN1(w0[3]), .IN2(n6), .Q(N16) );
  AND2X1 U16 ( .IN1(w0[2]), .IN2(n6), .Q(N15) );
  AND2X1 U17 ( .IN1(w0[1]), .IN2(n6), .Q(N14) );
  AND2X1 U18 ( .IN1(w0[0]), .IN2(n6), .Q(N13) );
  AND2X1 U19 ( .IN1(wrptr[8]), .IN2(n6), .Q(N12) );
  AND2X1 U20 ( .IN1(wrptr[7]), .IN2(n6), .Q(N11) );
  AND2X1 U21 ( .IN1(wrptr[6]), .IN2(n6), .Q(N10) );
  NOR2X0 U3 ( .IN1(n1), .IN2(flush), .QN(N19) );
  NOR2X0 U10 ( .IN1(n2), .IN2(flush), .QN(N20) );
  NOR2X0 U11 ( .IN1(n3), .IN2(flush), .QN(N21) );
  NBUFFX2 U12 ( .INP(rst), .Z(n4) );
  NBUFFX2 U22 ( .INP(rst), .Z(n5) );
  INVX0 U23 ( .INP(flush), .ZN(n6) );
endmodule


module flush_sync ( clk_in, rst, flush, sync_flush_BAR );
  input clk_in, rst, flush;
  output sync_flush_BAR;
  wire   f0;

  DFFARX1 f0_reg ( .D(flush), .CLK(clk_in), .RSTB(rst), .Q(f0) );
  DFFARX1 sync_flush_reg ( .D(f0), .CLK(clk_in), .RSTB(rst), .QN(
        sync_flush_BAR) );
endmodule


module memory_datasize32_addrbits8_depth128 ( clk_in, flush, rst, clk_out, 
        rden, rdaddr, wraddr, dataIn, dataOut, sync_flush_BAR, wren_BAR );
  input [7:0] rdaddr;
  input [7:0] wraddr;
  input [31:0] dataIn;
  output [31:0] dataOut;
  input clk_in, flush, rst, clk_out, rden, sync_flush_BAR, wren_BAR;
  wire   N15, N16, N17, N18, N19, N20, N21, sync_flush, wren, \FIFO[0][31] ,
         \FIFO[0][30] , \FIFO[0][29] , \FIFO[0][28] , \FIFO[0][27] ,
         \FIFO[0][26] , \FIFO[0][25] , \FIFO[0][24] , \FIFO[0][23] ,
         \FIFO[0][22] , \FIFO[0][21] , \FIFO[0][20] , \FIFO[0][19] ,
         \FIFO[0][18] , \FIFO[0][17] , \FIFO[0][16] , \FIFO[0][15] ,
         \FIFO[0][14] , \FIFO[0][13] , \FIFO[0][12] , \FIFO[0][11] ,
         \FIFO[0][10] , \FIFO[0][9] , \FIFO[0][8] , \FIFO[0][7] , \FIFO[0][6] ,
         \FIFO[0][5] , \FIFO[0][4] , \FIFO[0][3] , \FIFO[0][2] , \FIFO[0][1] ,
         \FIFO[0][0] , \FIFO[1][31] , \FIFO[1][30] , \FIFO[1][29] ,
         \FIFO[1][28] , \FIFO[1][27] , \FIFO[1][26] , \FIFO[1][25] ,
         \FIFO[1][24] , \FIFO[1][23] , \FIFO[1][22] , \FIFO[1][21] ,
         \FIFO[1][20] , \FIFO[1][19] , \FIFO[1][18] , \FIFO[1][17] ,
         \FIFO[1][16] , \FIFO[1][15] , \FIFO[1][14] , \FIFO[1][13] ,
         \FIFO[1][12] , \FIFO[1][11] , \FIFO[1][10] , \FIFO[1][9] ,
         \FIFO[1][8] , \FIFO[1][7] , \FIFO[1][6] , \FIFO[1][5] , \FIFO[1][4] ,
         \FIFO[1][3] , \FIFO[1][2] , \FIFO[1][1] , \FIFO[1][0] , \FIFO[2][31] ,
         \FIFO[2][30] , \FIFO[2][29] , \FIFO[2][28] , \FIFO[2][27] ,
         \FIFO[2][26] , \FIFO[2][25] , \FIFO[2][24] , \FIFO[2][23] ,
         \FIFO[2][22] , \FIFO[2][21] , \FIFO[2][20] , \FIFO[2][19] ,
         \FIFO[2][18] , \FIFO[2][17] , \FIFO[2][16] , \FIFO[2][15] ,
         \FIFO[2][14] , \FIFO[2][13] , \FIFO[2][12] , \FIFO[2][11] ,
         \FIFO[2][10] , \FIFO[2][9] , \FIFO[2][8] , \FIFO[2][7] , \FIFO[2][6] ,
         \FIFO[2][5] , \FIFO[2][4] , \FIFO[2][3] , \FIFO[2][2] , \FIFO[2][1] ,
         \FIFO[2][0] , \FIFO[3][31] , \FIFO[3][30] , \FIFO[3][29] ,
         \FIFO[3][28] , \FIFO[3][27] , \FIFO[3][26] , \FIFO[3][25] ,
         \FIFO[3][24] , \FIFO[3][23] , \FIFO[3][22] , \FIFO[3][21] ,
         \FIFO[3][20] , \FIFO[3][19] , \FIFO[3][18] , \FIFO[3][17] ,
         \FIFO[3][16] , \FIFO[3][15] , \FIFO[3][14] , \FIFO[3][13] ,
         \FIFO[3][12] , \FIFO[3][11] , \FIFO[3][10] , \FIFO[3][9] ,
         \FIFO[3][8] , \FIFO[3][7] , \FIFO[3][6] , \FIFO[3][5] , \FIFO[3][4] ,
         \FIFO[3][3] , \FIFO[3][2] , \FIFO[3][1] , \FIFO[3][0] , \FIFO[4][31] ,
         \FIFO[4][30] , \FIFO[4][29] , \FIFO[4][28] , \FIFO[4][27] ,
         \FIFO[4][26] , \FIFO[4][25] , \FIFO[4][24] , \FIFO[4][23] ,
         \FIFO[4][22] , \FIFO[4][21] , \FIFO[4][20] , \FIFO[4][19] ,
         \FIFO[4][18] , \FIFO[4][17] , \FIFO[4][16] , \FIFO[4][15] ,
         \FIFO[4][14] , \FIFO[4][13] , \FIFO[4][12] , \FIFO[4][11] ,
         \FIFO[4][10] , \FIFO[4][9] , \FIFO[4][8] , \FIFO[4][7] , \FIFO[4][6] ,
         \FIFO[4][5] , \FIFO[4][4] , \FIFO[4][3] , \FIFO[4][2] , \FIFO[4][1] ,
         \FIFO[4][0] , \FIFO[5][31] , \FIFO[5][30] , \FIFO[5][29] ,
         \FIFO[5][28] , \FIFO[5][27] , \FIFO[5][26] , \FIFO[5][25] ,
         \FIFO[5][24] , \FIFO[5][23] , \FIFO[5][22] , \FIFO[5][21] ,
         \FIFO[5][20] , \FIFO[5][19] , \FIFO[5][18] , \FIFO[5][17] ,
         \FIFO[5][16] , \FIFO[5][15] , \FIFO[5][14] , \FIFO[5][13] ,
         \FIFO[5][12] , \FIFO[5][11] , \FIFO[5][10] , \FIFO[5][9] ,
         \FIFO[5][8] , \FIFO[5][7] , \FIFO[5][6] , \FIFO[5][5] , \FIFO[5][4] ,
         \FIFO[5][3] , \FIFO[5][2] , \FIFO[5][1] , \FIFO[5][0] , \FIFO[6][31] ,
         \FIFO[6][30] , \FIFO[6][29] , \FIFO[6][28] , \FIFO[6][27] ,
         \FIFO[6][26] , \FIFO[6][25] , \FIFO[6][24] , \FIFO[6][23] ,
         \FIFO[6][22] , \FIFO[6][21] , \FIFO[6][20] , \FIFO[6][19] ,
         \FIFO[6][18] , \FIFO[6][17] , \FIFO[6][16] , \FIFO[6][15] ,
         \FIFO[6][14] , \FIFO[6][13] , \FIFO[6][12] , \FIFO[6][11] ,
         \FIFO[6][10] , \FIFO[6][9] , \FIFO[6][8] , \FIFO[6][7] , \FIFO[6][6] ,
         \FIFO[6][5] , \FIFO[6][4] , \FIFO[6][3] , \FIFO[6][2] , \FIFO[6][1] ,
         \FIFO[6][0] , \FIFO[7][31] , \FIFO[7][30] , \FIFO[7][29] ,
         \FIFO[7][28] , \FIFO[7][27] , \FIFO[7][26] , \FIFO[7][25] ,
         \FIFO[7][24] , \FIFO[7][23] , \FIFO[7][22] , \FIFO[7][21] ,
         \FIFO[7][20] , \FIFO[7][19] , \FIFO[7][18] , \FIFO[7][17] ,
         \FIFO[7][16] , \FIFO[7][15] , \FIFO[7][14] , \FIFO[7][13] ,
         \FIFO[7][12] , \FIFO[7][11] , \FIFO[7][10] , \FIFO[7][9] ,
         \FIFO[7][8] , \FIFO[7][7] , \FIFO[7][6] , \FIFO[7][5] , \FIFO[7][4] ,
         \FIFO[7][3] , \FIFO[7][2] , \FIFO[7][1] , \FIFO[7][0] , \FIFO[8][31] ,
         \FIFO[8][30] , \FIFO[8][29] , \FIFO[8][28] , \FIFO[8][27] ,
         \FIFO[8][26] , \FIFO[8][25] , \FIFO[8][24] , \FIFO[8][23] ,
         \FIFO[8][22] , \FIFO[8][21] , \FIFO[8][20] , \FIFO[8][19] ,
         \FIFO[8][18] , \FIFO[8][17] , \FIFO[8][16] , \FIFO[8][15] ,
         \FIFO[8][14] , \FIFO[8][13] , \FIFO[8][12] , \FIFO[8][11] ,
         \FIFO[8][10] , \FIFO[8][9] , \FIFO[8][8] , \FIFO[8][7] , \FIFO[8][6] ,
         \FIFO[8][5] , \FIFO[8][4] , \FIFO[8][3] , \FIFO[8][2] , \FIFO[8][1] ,
         \FIFO[8][0] , \FIFO[9][31] , \FIFO[9][30] , \FIFO[9][29] ,
         \FIFO[9][28] , \FIFO[9][27] , \FIFO[9][26] , \FIFO[9][25] ,
         \FIFO[9][24] , \FIFO[9][23] , \FIFO[9][22] , \FIFO[9][21] ,
         \FIFO[9][20] , \FIFO[9][19] , \FIFO[9][18] , \FIFO[9][17] ,
         \FIFO[9][16] , \FIFO[9][15] , \FIFO[9][14] , \FIFO[9][13] ,
         \FIFO[9][12] , \FIFO[9][11] , \FIFO[9][10] , \FIFO[9][9] ,
         \FIFO[9][8] , \FIFO[9][7] , \FIFO[9][6] , \FIFO[9][5] , \FIFO[9][4] ,
         \FIFO[9][3] , \FIFO[9][2] , \FIFO[9][1] , \FIFO[9][0] ,
         \FIFO[10][31] , \FIFO[10][30] , \FIFO[10][29] , \FIFO[10][28] ,
         \FIFO[10][27] , \FIFO[10][26] , \FIFO[10][25] , \FIFO[10][24] ,
         \FIFO[10][23] , \FIFO[10][22] , \FIFO[10][21] , \FIFO[10][20] ,
         \FIFO[10][19] , \FIFO[10][18] , \FIFO[10][17] , \FIFO[10][16] ,
         \FIFO[10][15] , \FIFO[10][14] , \FIFO[10][13] , \FIFO[10][12] ,
         \FIFO[10][11] , \FIFO[10][10] , \FIFO[10][9] , \FIFO[10][8] ,
         \FIFO[10][7] , \FIFO[10][6] , \FIFO[10][5] , \FIFO[10][4] ,
         \FIFO[10][3] , \FIFO[10][2] , \FIFO[10][1] , \FIFO[10][0] ,
         \FIFO[11][31] , \FIFO[11][30] , \FIFO[11][29] , \FIFO[11][28] ,
         \FIFO[11][27] , \FIFO[11][26] , \FIFO[11][25] , \FIFO[11][24] ,
         \FIFO[11][23] , \FIFO[11][22] , \FIFO[11][21] , \FIFO[11][20] ,
         \FIFO[11][19] , \FIFO[11][18] , \FIFO[11][17] , \FIFO[11][16] ,
         \FIFO[11][15] , \FIFO[11][14] , \FIFO[11][13] , \FIFO[11][12] ,
         \FIFO[11][11] , \FIFO[11][10] , \FIFO[11][9] , \FIFO[11][8] ,
         \FIFO[11][7] , \FIFO[11][6] , \FIFO[11][5] , \FIFO[11][4] ,
         \FIFO[11][3] , \FIFO[11][2] , \FIFO[11][1] , \FIFO[11][0] ,
         \FIFO[12][31] , \FIFO[12][30] , \FIFO[12][29] , \FIFO[12][28] ,
         \FIFO[12][27] , \FIFO[12][26] , \FIFO[12][25] , \FIFO[12][24] ,
         \FIFO[12][23] , \FIFO[12][22] , \FIFO[12][21] , \FIFO[12][20] ,
         \FIFO[12][19] , \FIFO[12][18] , \FIFO[12][17] , \FIFO[12][16] ,
         \FIFO[12][15] , \FIFO[12][14] , \FIFO[12][13] , \FIFO[12][12] ,
         \FIFO[12][11] , \FIFO[12][10] , \FIFO[12][9] , \FIFO[12][8] ,
         \FIFO[12][7] , \FIFO[12][6] , \FIFO[12][5] , \FIFO[12][4] ,
         \FIFO[12][3] , \FIFO[12][2] , \FIFO[12][1] , \FIFO[12][0] ,
         \FIFO[13][31] , \FIFO[13][30] , \FIFO[13][29] , \FIFO[13][28] ,
         \FIFO[13][27] , \FIFO[13][26] , \FIFO[13][25] , \FIFO[13][24] ,
         \FIFO[13][23] , \FIFO[13][22] , \FIFO[13][21] , \FIFO[13][20] ,
         \FIFO[13][19] , \FIFO[13][18] , \FIFO[13][17] , \FIFO[13][16] ,
         \FIFO[13][15] , \FIFO[13][14] , \FIFO[13][13] , \FIFO[13][12] ,
         \FIFO[13][11] , \FIFO[13][10] , \FIFO[13][9] , \FIFO[13][8] ,
         \FIFO[13][7] , \FIFO[13][6] , \FIFO[13][5] , \FIFO[13][4] ,
         \FIFO[13][3] , \FIFO[13][2] , \FIFO[13][1] , \FIFO[13][0] ,
         \FIFO[14][31] , \FIFO[14][30] , \FIFO[14][29] , \FIFO[14][28] ,
         \FIFO[14][27] , \FIFO[14][26] , \FIFO[14][25] , \FIFO[14][24] ,
         \FIFO[14][23] , \FIFO[14][22] , \FIFO[14][21] , \FIFO[14][20] ,
         \FIFO[14][19] , \FIFO[14][18] , \FIFO[14][17] , \FIFO[14][16] ,
         \FIFO[14][15] , \FIFO[14][14] , \FIFO[14][13] , \FIFO[14][12] ,
         \FIFO[14][11] , \FIFO[14][10] , \FIFO[14][9] , \FIFO[14][8] ,
         \FIFO[14][7] , \FIFO[14][6] , \FIFO[14][5] , \FIFO[14][4] ,
         \FIFO[14][3] , \FIFO[14][2] , \FIFO[14][1] , \FIFO[14][0] ,
         \FIFO[15][31] , \FIFO[15][30] , \FIFO[15][29] , \FIFO[15][28] ,
         \FIFO[15][27] , \FIFO[15][26] , \FIFO[15][25] , \FIFO[15][24] ,
         \FIFO[15][23] , \FIFO[15][22] , \FIFO[15][21] , \FIFO[15][20] ,
         \FIFO[15][19] , \FIFO[15][18] , \FIFO[15][17] , \FIFO[15][16] ,
         \FIFO[15][15] , \FIFO[15][14] , \FIFO[15][13] , \FIFO[15][12] ,
         \FIFO[15][11] , \FIFO[15][10] , \FIFO[15][9] , \FIFO[15][8] ,
         \FIFO[15][7] , \FIFO[15][6] , \FIFO[15][5] , \FIFO[15][4] ,
         \FIFO[15][3] , \FIFO[15][2] , \FIFO[15][1] , \FIFO[15][0] ,
         \FIFO[16][31] , \FIFO[16][30] , \FIFO[16][29] , \FIFO[16][28] ,
         \FIFO[16][27] , \FIFO[16][26] , \FIFO[16][25] , \FIFO[16][24] ,
         \FIFO[16][23] , \FIFO[16][22] , \FIFO[16][21] , \FIFO[16][20] ,
         \FIFO[16][19] , \FIFO[16][18] , \FIFO[16][17] , \FIFO[16][16] ,
         \FIFO[16][15] , \FIFO[16][14] , \FIFO[16][13] , \FIFO[16][12] ,
         \FIFO[16][11] , \FIFO[16][10] , \FIFO[16][9] , \FIFO[16][8] ,
         \FIFO[16][7] , \FIFO[16][6] , \FIFO[16][5] , \FIFO[16][4] ,
         \FIFO[16][3] , \FIFO[16][2] , \FIFO[16][1] , \FIFO[16][0] ,
         \FIFO[17][31] , \FIFO[17][30] , \FIFO[17][29] , \FIFO[17][28] ,
         \FIFO[17][27] , \FIFO[17][26] , \FIFO[17][25] , \FIFO[17][24] ,
         \FIFO[17][23] , \FIFO[17][22] , \FIFO[17][21] , \FIFO[17][20] ,
         \FIFO[17][19] , \FIFO[17][18] , \FIFO[17][17] , \FIFO[17][16] ,
         \FIFO[17][15] , \FIFO[17][14] , \FIFO[17][13] , \FIFO[17][12] ,
         \FIFO[17][11] , \FIFO[17][10] , \FIFO[17][9] , \FIFO[17][8] ,
         \FIFO[17][7] , \FIFO[17][6] , \FIFO[17][5] , \FIFO[17][4] ,
         \FIFO[17][3] , \FIFO[17][2] , \FIFO[17][1] , \FIFO[17][0] ,
         \FIFO[18][31] , \FIFO[18][30] , \FIFO[18][29] , \FIFO[18][28] ,
         \FIFO[18][27] , \FIFO[18][26] , \FIFO[18][25] , \FIFO[18][24] ,
         \FIFO[18][23] , \FIFO[18][22] , \FIFO[18][21] , \FIFO[18][20] ,
         \FIFO[18][19] , \FIFO[18][18] , \FIFO[18][17] , \FIFO[18][16] ,
         \FIFO[18][15] , \FIFO[18][14] , \FIFO[18][13] , \FIFO[18][12] ,
         \FIFO[18][11] , \FIFO[18][10] , \FIFO[18][9] , \FIFO[18][8] ,
         \FIFO[18][7] , \FIFO[18][6] , \FIFO[18][5] , \FIFO[18][4] ,
         \FIFO[18][3] , \FIFO[18][2] , \FIFO[18][1] , \FIFO[18][0] ,
         \FIFO[19][31] , \FIFO[19][30] , \FIFO[19][29] , \FIFO[19][28] ,
         \FIFO[19][27] , \FIFO[19][26] , \FIFO[19][25] , \FIFO[19][24] ,
         \FIFO[19][23] , \FIFO[19][22] , \FIFO[19][21] , \FIFO[19][20] ,
         \FIFO[19][19] , \FIFO[19][18] , \FIFO[19][17] , \FIFO[19][16] ,
         \FIFO[19][15] , \FIFO[19][14] , \FIFO[19][13] , \FIFO[19][12] ,
         \FIFO[19][11] , \FIFO[19][10] , \FIFO[19][9] , \FIFO[19][8] ,
         \FIFO[19][7] , \FIFO[19][6] , \FIFO[19][5] , \FIFO[19][4] ,
         \FIFO[19][3] , \FIFO[19][2] , \FIFO[19][1] , \FIFO[19][0] ,
         \FIFO[20][31] , \FIFO[20][30] , \FIFO[20][29] , \FIFO[20][28] ,
         \FIFO[20][27] , \FIFO[20][26] , \FIFO[20][25] , \FIFO[20][24] ,
         \FIFO[20][23] , \FIFO[20][22] , \FIFO[20][21] , \FIFO[20][20] ,
         \FIFO[20][19] , \FIFO[20][18] , \FIFO[20][17] , \FIFO[20][16] ,
         \FIFO[20][15] , \FIFO[20][14] , \FIFO[20][13] , \FIFO[20][12] ,
         \FIFO[20][11] , \FIFO[20][10] , \FIFO[20][9] , \FIFO[20][8] ,
         \FIFO[20][7] , \FIFO[20][6] , \FIFO[20][5] , \FIFO[20][4] ,
         \FIFO[20][3] , \FIFO[20][2] , \FIFO[20][1] , \FIFO[20][0] ,
         \FIFO[21][31] , \FIFO[21][30] , \FIFO[21][29] , \FIFO[21][28] ,
         \FIFO[21][27] , \FIFO[21][26] , \FIFO[21][25] , \FIFO[21][24] ,
         \FIFO[21][23] , \FIFO[21][22] , \FIFO[21][21] , \FIFO[21][20] ,
         \FIFO[21][19] , \FIFO[21][18] , \FIFO[21][17] , \FIFO[21][16] ,
         \FIFO[21][15] , \FIFO[21][14] , \FIFO[21][13] , \FIFO[21][12] ,
         \FIFO[21][11] , \FIFO[21][10] , \FIFO[21][9] , \FIFO[21][8] ,
         \FIFO[21][7] , \FIFO[21][6] , \FIFO[21][5] , \FIFO[21][4] ,
         \FIFO[21][3] , \FIFO[21][2] , \FIFO[21][1] , \FIFO[21][0] ,
         \FIFO[22][31] , \FIFO[22][30] , \FIFO[22][29] , \FIFO[22][28] ,
         \FIFO[22][27] , \FIFO[22][26] , \FIFO[22][25] , \FIFO[22][24] ,
         \FIFO[22][23] , \FIFO[22][22] , \FIFO[22][21] , \FIFO[22][20] ,
         \FIFO[22][19] , \FIFO[22][18] , \FIFO[22][17] , \FIFO[22][16] ,
         \FIFO[22][15] , \FIFO[22][14] , \FIFO[22][13] , \FIFO[22][12] ,
         \FIFO[22][11] , \FIFO[22][10] , \FIFO[22][9] , \FIFO[22][8] ,
         \FIFO[22][7] , \FIFO[22][6] , \FIFO[22][5] , \FIFO[22][4] ,
         \FIFO[22][3] , \FIFO[22][2] , \FIFO[22][1] , \FIFO[22][0] ,
         \FIFO[23][31] , \FIFO[23][30] , \FIFO[23][29] , \FIFO[23][28] ,
         \FIFO[23][27] , \FIFO[23][26] , \FIFO[23][25] , \FIFO[23][24] ,
         \FIFO[23][23] , \FIFO[23][22] , \FIFO[23][21] , \FIFO[23][20] ,
         \FIFO[23][19] , \FIFO[23][18] , \FIFO[23][17] , \FIFO[23][16] ,
         \FIFO[23][15] , \FIFO[23][14] , \FIFO[23][13] , \FIFO[23][12] ,
         \FIFO[23][11] , \FIFO[23][10] , \FIFO[23][9] , \FIFO[23][8] ,
         \FIFO[23][7] , \FIFO[23][6] , \FIFO[23][5] , \FIFO[23][4] ,
         \FIFO[23][3] , \FIFO[23][2] , \FIFO[23][1] , \FIFO[23][0] ,
         \FIFO[24][31] , \FIFO[24][30] , \FIFO[24][29] , \FIFO[24][28] ,
         \FIFO[24][27] , \FIFO[24][26] , \FIFO[24][25] , \FIFO[24][24] ,
         \FIFO[24][23] , \FIFO[24][22] , \FIFO[24][21] , \FIFO[24][20] ,
         \FIFO[24][19] , \FIFO[24][18] , \FIFO[24][17] , \FIFO[24][16] ,
         \FIFO[24][15] , \FIFO[24][14] , \FIFO[24][13] , \FIFO[24][12] ,
         \FIFO[24][11] , \FIFO[24][10] , \FIFO[24][9] , \FIFO[24][8] ,
         \FIFO[24][7] , \FIFO[24][6] , \FIFO[24][5] , \FIFO[24][4] ,
         \FIFO[24][3] , \FIFO[24][2] , \FIFO[24][1] , \FIFO[24][0] ,
         \FIFO[25][31] , \FIFO[25][30] , \FIFO[25][29] , \FIFO[25][28] ,
         \FIFO[25][27] , \FIFO[25][26] , \FIFO[25][25] , \FIFO[25][24] ,
         \FIFO[25][23] , \FIFO[25][22] , \FIFO[25][21] , \FIFO[25][20] ,
         \FIFO[25][19] , \FIFO[25][18] , \FIFO[25][17] , \FIFO[25][16] ,
         \FIFO[25][15] , \FIFO[25][14] , \FIFO[25][13] , \FIFO[25][12] ,
         \FIFO[25][11] , \FIFO[25][10] , \FIFO[25][9] , \FIFO[25][8] ,
         \FIFO[25][7] , \FIFO[25][6] , \FIFO[25][5] , \FIFO[25][4] ,
         \FIFO[25][3] , \FIFO[25][2] , \FIFO[25][1] , \FIFO[25][0] ,
         \FIFO[26][31] , \FIFO[26][30] , \FIFO[26][29] , \FIFO[26][28] ,
         \FIFO[26][27] , \FIFO[26][26] , \FIFO[26][25] , \FIFO[26][24] ,
         \FIFO[26][23] , \FIFO[26][22] , \FIFO[26][21] , \FIFO[26][20] ,
         \FIFO[26][19] , \FIFO[26][18] , \FIFO[26][17] , \FIFO[26][16] ,
         \FIFO[26][15] , \FIFO[26][14] , \FIFO[26][13] , \FIFO[26][12] ,
         \FIFO[26][11] , \FIFO[26][10] , \FIFO[26][9] , \FIFO[26][8] ,
         \FIFO[26][7] , \FIFO[26][6] , \FIFO[26][5] , \FIFO[26][4] ,
         \FIFO[26][3] , \FIFO[26][2] , \FIFO[26][1] , \FIFO[26][0] ,
         \FIFO[27][31] , \FIFO[27][30] , \FIFO[27][29] , \FIFO[27][28] ,
         \FIFO[27][27] , \FIFO[27][26] , \FIFO[27][25] , \FIFO[27][24] ,
         \FIFO[27][23] , \FIFO[27][22] , \FIFO[27][21] , \FIFO[27][20] ,
         \FIFO[27][19] , \FIFO[27][18] , \FIFO[27][17] , \FIFO[27][16] ,
         \FIFO[27][15] , \FIFO[27][14] , \FIFO[27][13] , \FIFO[27][12] ,
         \FIFO[27][11] , \FIFO[27][10] , \FIFO[27][9] , \FIFO[27][8] ,
         \FIFO[27][7] , \FIFO[27][6] , \FIFO[27][5] , \FIFO[27][4] ,
         \FIFO[27][3] , \FIFO[27][2] , \FIFO[27][1] , \FIFO[27][0] ,
         \FIFO[28][31] , \FIFO[28][30] , \FIFO[28][29] , \FIFO[28][28] ,
         \FIFO[28][27] , \FIFO[28][26] , \FIFO[28][25] , \FIFO[28][24] ,
         \FIFO[28][23] , \FIFO[28][22] , \FIFO[28][21] , \FIFO[28][20] ,
         \FIFO[28][19] , \FIFO[28][18] , \FIFO[28][17] , \FIFO[28][16] ,
         \FIFO[28][15] , \FIFO[28][14] , \FIFO[28][13] , \FIFO[28][12] ,
         \FIFO[28][11] , \FIFO[28][10] , \FIFO[28][9] , \FIFO[28][8] ,
         \FIFO[28][7] , \FIFO[28][6] , \FIFO[28][5] , \FIFO[28][4] ,
         \FIFO[28][3] , \FIFO[28][2] , \FIFO[28][1] , \FIFO[28][0] ,
         \FIFO[29][31] , \FIFO[29][30] , \FIFO[29][29] , \FIFO[29][28] ,
         \FIFO[29][27] , \FIFO[29][26] , \FIFO[29][25] , \FIFO[29][24] ,
         \FIFO[29][23] , \FIFO[29][22] , \FIFO[29][21] , \FIFO[29][20] ,
         \FIFO[29][19] , \FIFO[29][18] , \FIFO[29][17] , \FIFO[29][16] ,
         \FIFO[29][15] , \FIFO[29][14] , \FIFO[29][13] , \FIFO[29][12] ,
         \FIFO[29][11] , \FIFO[29][10] , \FIFO[29][9] , \FIFO[29][8] ,
         \FIFO[29][7] , \FIFO[29][6] , \FIFO[29][5] , \FIFO[29][4] ,
         \FIFO[29][3] , \FIFO[29][2] , \FIFO[29][1] , \FIFO[29][0] ,
         \FIFO[30][31] , \FIFO[30][30] , \FIFO[30][29] , \FIFO[30][28] ,
         \FIFO[30][27] , \FIFO[30][26] , \FIFO[30][25] , \FIFO[30][24] ,
         \FIFO[30][23] , \FIFO[30][22] , \FIFO[30][21] , \FIFO[30][20] ,
         \FIFO[30][19] , \FIFO[30][18] , \FIFO[30][17] , \FIFO[30][16] ,
         \FIFO[30][15] , \FIFO[30][14] , \FIFO[30][13] , \FIFO[30][12] ,
         \FIFO[30][11] , \FIFO[30][10] , \FIFO[30][9] , \FIFO[30][8] ,
         \FIFO[30][7] , \FIFO[30][6] , \FIFO[30][5] , \FIFO[30][4] ,
         \FIFO[30][3] , \FIFO[30][2] , \FIFO[30][1] , \FIFO[30][0] ,
         \FIFO[31][31] , \FIFO[31][30] , \FIFO[31][29] , \FIFO[31][28] ,
         \FIFO[31][27] , \FIFO[31][26] , \FIFO[31][25] , \FIFO[31][24] ,
         \FIFO[31][23] , \FIFO[31][22] , \FIFO[31][21] , \FIFO[31][20] ,
         \FIFO[31][19] , \FIFO[31][18] , \FIFO[31][17] , \FIFO[31][16] ,
         \FIFO[31][15] , \FIFO[31][14] , \FIFO[31][13] , \FIFO[31][12] ,
         \FIFO[31][11] , \FIFO[31][10] , \FIFO[31][9] , \FIFO[31][8] ,
         \FIFO[31][7] , \FIFO[31][6] , \FIFO[31][5] , \FIFO[31][4] ,
         \FIFO[31][3] , \FIFO[31][2] , \FIFO[31][1] , \FIFO[31][0] ,
         \FIFO[32][31] , \FIFO[32][30] , \FIFO[32][29] , \FIFO[32][28] ,
         \FIFO[32][27] , \FIFO[32][26] , \FIFO[32][25] , \FIFO[32][24] ,
         \FIFO[32][23] , \FIFO[32][22] , \FIFO[32][21] , \FIFO[32][20] ,
         \FIFO[32][19] , \FIFO[32][18] , \FIFO[32][17] , \FIFO[32][16] ,
         \FIFO[32][15] , \FIFO[32][14] , \FIFO[32][13] , \FIFO[32][12] ,
         \FIFO[32][11] , \FIFO[32][10] , \FIFO[32][9] , \FIFO[32][8] ,
         \FIFO[32][7] , \FIFO[32][6] , \FIFO[32][5] , \FIFO[32][4] ,
         \FIFO[32][3] , \FIFO[32][2] , \FIFO[32][1] , \FIFO[32][0] ,
         \FIFO[33][31] , \FIFO[33][30] , \FIFO[33][29] , \FIFO[33][28] ,
         \FIFO[33][27] , \FIFO[33][26] , \FIFO[33][25] , \FIFO[33][24] ,
         \FIFO[33][23] , \FIFO[33][22] , \FIFO[33][21] , \FIFO[33][20] ,
         \FIFO[33][19] , \FIFO[33][18] , \FIFO[33][17] , \FIFO[33][16] ,
         \FIFO[33][15] , \FIFO[33][14] , \FIFO[33][13] , \FIFO[33][12] ,
         \FIFO[33][11] , \FIFO[33][10] , \FIFO[33][9] , \FIFO[33][8] ,
         \FIFO[33][7] , \FIFO[33][6] , \FIFO[33][5] , \FIFO[33][4] ,
         \FIFO[33][3] , \FIFO[33][2] , \FIFO[33][1] , \FIFO[33][0] ,
         \FIFO[34][31] , \FIFO[34][30] , \FIFO[34][29] , \FIFO[34][28] ,
         \FIFO[34][27] , \FIFO[34][26] , \FIFO[34][25] , \FIFO[34][24] ,
         \FIFO[34][23] , \FIFO[34][22] , \FIFO[34][21] , \FIFO[34][20] ,
         \FIFO[34][19] , \FIFO[34][18] , \FIFO[34][17] , \FIFO[34][16] ,
         \FIFO[34][15] , \FIFO[34][14] , \FIFO[34][13] , \FIFO[34][12] ,
         \FIFO[34][11] , \FIFO[34][10] , \FIFO[34][9] , \FIFO[34][8] ,
         \FIFO[34][7] , \FIFO[34][6] , \FIFO[34][5] , \FIFO[34][4] ,
         \FIFO[34][3] , \FIFO[34][2] , \FIFO[34][1] , \FIFO[34][0] ,
         \FIFO[35][31] , \FIFO[35][30] , \FIFO[35][29] , \FIFO[35][28] ,
         \FIFO[35][27] , \FIFO[35][26] , \FIFO[35][25] , \FIFO[35][24] ,
         \FIFO[35][23] , \FIFO[35][22] , \FIFO[35][21] , \FIFO[35][20] ,
         \FIFO[35][19] , \FIFO[35][18] , \FIFO[35][17] , \FIFO[35][16] ,
         \FIFO[35][15] , \FIFO[35][14] , \FIFO[35][13] , \FIFO[35][12] ,
         \FIFO[35][11] , \FIFO[35][10] , \FIFO[35][9] , \FIFO[35][8] ,
         \FIFO[35][7] , \FIFO[35][6] , \FIFO[35][5] , \FIFO[35][4] ,
         \FIFO[35][3] , \FIFO[35][2] , \FIFO[35][1] , \FIFO[35][0] ,
         \FIFO[36][31] , \FIFO[36][30] , \FIFO[36][29] , \FIFO[36][28] ,
         \FIFO[36][27] , \FIFO[36][26] , \FIFO[36][25] , \FIFO[36][24] ,
         \FIFO[36][23] , \FIFO[36][22] , \FIFO[36][21] , \FIFO[36][20] ,
         \FIFO[36][19] , \FIFO[36][18] , \FIFO[36][17] , \FIFO[36][16] ,
         \FIFO[36][15] , \FIFO[36][14] , \FIFO[36][13] , \FIFO[36][12] ,
         \FIFO[36][11] , \FIFO[36][10] , \FIFO[36][9] , \FIFO[36][8] ,
         \FIFO[36][7] , \FIFO[36][6] , \FIFO[36][5] , \FIFO[36][4] ,
         \FIFO[36][3] , \FIFO[36][2] , \FIFO[36][1] , \FIFO[36][0] ,
         \FIFO[37][31] , \FIFO[37][30] , \FIFO[37][29] , \FIFO[37][28] ,
         \FIFO[37][27] , \FIFO[37][26] , \FIFO[37][25] , \FIFO[37][24] ,
         \FIFO[37][23] , \FIFO[37][22] , \FIFO[37][21] , \FIFO[37][20] ,
         \FIFO[37][19] , \FIFO[37][18] , \FIFO[37][17] , \FIFO[37][16] ,
         \FIFO[37][15] , \FIFO[37][14] , \FIFO[37][13] , \FIFO[37][12] ,
         \FIFO[37][11] , \FIFO[37][10] , \FIFO[37][9] , \FIFO[37][8] ,
         \FIFO[37][7] , \FIFO[37][6] , \FIFO[37][5] , \FIFO[37][4] ,
         \FIFO[37][3] , \FIFO[37][2] , \FIFO[37][1] , \FIFO[37][0] ,
         \FIFO[38][31] , \FIFO[38][30] , \FIFO[38][29] , \FIFO[38][28] ,
         \FIFO[38][27] , \FIFO[38][26] , \FIFO[38][25] , \FIFO[38][24] ,
         \FIFO[38][23] , \FIFO[38][22] , \FIFO[38][21] , \FIFO[38][20] ,
         \FIFO[38][19] , \FIFO[38][18] , \FIFO[38][17] , \FIFO[38][16] ,
         \FIFO[38][15] , \FIFO[38][14] , \FIFO[38][13] , \FIFO[38][12] ,
         \FIFO[38][11] , \FIFO[38][10] , \FIFO[38][9] , \FIFO[38][8] ,
         \FIFO[38][7] , \FIFO[38][6] , \FIFO[38][5] , \FIFO[38][4] ,
         \FIFO[38][3] , \FIFO[38][2] , \FIFO[38][1] , \FIFO[38][0] ,
         \FIFO[39][31] , \FIFO[39][30] , \FIFO[39][29] , \FIFO[39][28] ,
         \FIFO[39][27] , \FIFO[39][26] , \FIFO[39][25] , \FIFO[39][24] ,
         \FIFO[39][23] , \FIFO[39][22] , \FIFO[39][21] , \FIFO[39][20] ,
         \FIFO[39][19] , \FIFO[39][18] , \FIFO[39][17] , \FIFO[39][16] ,
         \FIFO[39][15] , \FIFO[39][14] , \FIFO[39][13] , \FIFO[39][12] ,
         \FIFO[39][11] , \FIFO[39][10] , \FIFO[39][9] , \FIFO[39][8] ,
         \FIFO[39][7] , \FIFO[39][6] , \FIFO[39][5] , \FIFO[39][4] ,
         \FIFO[39][3] , \FIFO[39][2] , \FIFO[39][1] , \FIFO[39][0] ,
         \FIFO[40][31] , \FIFO[40][30] , \FIFO[40][29] , \FIFO[40][28] ,
         \FIFO[40][27] , \FIFO[40][26] , \FIFO[40][25] , \FIFO[40][24] ,
         \FIFO[40][23] , \FIFO[40][22] , \FIFO[40][21] , \FIFO[40][20] ,
         \FIFO[40][19] , \FIFO[40][18] , \FIFO[40][17] , \FIFO[40][16] ,
         \FIFO[40][15] , \FIFO[40][14] , \FIFO[40][13] , \FIFO[40][12] ,
         \FIFO[40][11] , \FIFO[40][10] , \FIFO[40][9] , \FIFO[40][8] ,
         \FIFO[40][7] , \FIFO[40][6] , \FIFO[40][5] , \FIFO[40][4] ,
         \FIFO[40][3] , \FIFO[40][2] , \FIFO[40][1] , \FIFO[40][0] ,
         \FIFO[41][31] , \FIFO[41][30] , \FIFO[41][29] , \FIFO[41][28] ,
         \FIFO[41][27] , \FIFO[41][26] , \FIFO[41][25] , \FIFO[41][24] ,
         \FIFO[41][23] , \FIFO[41][22] , \FIFO[41][21] , \FIFO[41][20] ,
         \FIFO[41][19] , \FIFO[41][18] , \FIFO[41][17] , \FIFO[41][16] ,
         \FIFO[41][15] , \FIFO[41][14] , \FIFO[41][13] , \FIFO[41][12] ,
         \FIFO[41][11] , \FIFO[41][10] , \FIFO[41][9] , \FIFO[41][8] ,
         \FIFO[41][7] , \FIFO[41][6] , \FIFO[41][5] , \FIFO[41][4] ,
         \FIFO[41][3] , \FIFO[41][2] , \FIFO[41][1] , \FIFO[41][0] ,
         \FIFO[42][31] , \FIFO[42][30] , \FIFO[42][29] , \FIFO[42][28] ,
         \FIFO[42][27] , \FIFO[42][26] , \FIFO[42][25] , \FIFO[42][24] ,
         \FIFO[42][23] , \FIFO[42][22] , \FIFO[42][21] , \FIFO[42][20] ,
         \FIFO[42][19] , \FIFO[42][18] , \FIFO[42][17] , \FIFO[42][16] ,
         \FIFO[42][15] , \FIFO[42][14] , \FIFO[42][13] , \FIFO[42][12] ,
         \FIFO[42][11] , \FIFO[42][10] , \FIFO[42][9] , \FIFO[42][8] ,
         \FIFO[42][7] , \FIFO[42][6] , \FIFO[42][5] , \FIFO[42][4] ,
         \FIFO[42][3] , \FIFO[42][2] , \FIFO[42][1] , \FIFO[42][0] ,
         \FIFO[43][31] , \FIFO[43][30] , \FIFO[43][29] , \FIFO[43][28] ,
         \FIFO[43][27] , \FIFO[43][26] , \FIFO[43][25] , \FIFO[43][24] ,
         \FIFO[43][23] , \FIFO[43][22] , \FIFO[43][21] , \FIFO[43][20] ,
         \FIFO[43][19] , \FIFO[43][18] , \FIFO[43][17] , \FIFO[43][16] ,
         \FIFO[43][15] , \FIFO[43][14] , \FIFO[43][13] , \FIFO[43][12] ,
         \FIFO[43][11] , \FIFO[43][10] , \FIFO[43][9] , \FIFO[43][8] ,
         \FIFO[43][7] , \FIFO[43][6] , \FIFO[43][5] , \FIFO[43][4] ,
         \FIFO[43][3] , \FIFO[43][2] , \FIFO[43][1] , \FIFO[43][0] ,
         \FIFO[44][31] , \FIFO[44][30] , \FIFO[44][29] , \FIFO[44][28] ,
         \FIFO[44][27] , \FIFO[44][26] , \FIFO[44][25] , \FIFO[44][24] ,
         \FIFO[44][23] , \FIFO[44][22] , \FIFO[44][21] , \FIFO[44][20] ,
         \FIFO[44][19] , \FIFO[44][18] , \FIFO[44][17] , \FIFO[44][16] ,
         \FIFO[44][15] , \FIFO[44][14] , \FIFO[44][13] , \FIFO[44][12] ,
         \FIFO[44][11] , \FIFO[44][10] , \FIFO[44][9] , \FIFO[44][8] ,
         \FIFO[44][7] , \FIFO[44][6] , \FIFO[44][5] , \FIFO[44][4] ,
         \FIFO[44][3] , \FIFO[44][2] , \FIFO[44][1] , \FIFO[44][0] ,
         \FIFO[45][31] , \FIFO[45][30] , \FIFO[45][29] , \FIFO[45][28] ,
         \FIFO[45][27] , \FIFO[45][26] , \FIFO[45][25] , \FIFO[45][24] ,
         \FIFO[45][23] , \FIFO[45][22] , \FIFO[45][21] , \FIFO[45][20] ,
         \FIFO[45][19] , \FIFO[45][18] , \FIFO[45][17] , \FIFO[45][16] ,
         \FIFO[45][15] , \FIFO[45][14] , \FIFO[45][13] , \FIFO[45][12] ,
         \FIFO[45][11] , \FIFO[45][10] , \FIFO[45][9] , \FIFO[45][8] ,
         \FIFO[45][7] , \FIFO[45][6] , \FIFO[45][5] , \FIFO[45][4] ,
         \FIFO[45][3] , \FIFO[45][2] , \FIFO[45][1] , \FIFO[45][0] ,
         \FIFO[46][31] , \FIFO[46][30] , \FIFO[46][29] , \FIFO[46][28] ,
         \FIFO[46][27] , \FIFO[46][26] , \FIFO[46][25] , \FIFO[46][24] ,
         \FIFO[46][23] , \FIFO[46][22] , \FIFO[46][21] , \FIFO[46][20] ,
         \FIFO[46][19] , \FIFO[46][18] , \FIFO[46][17] , \FIFO[46][16] ,
         \FIFO[46][15] , \FIFO[46][14] , \FIFO[46][13] , \FIFO[46][12] ,
         \FIFO[46][11] , \FIFO[46][10] , \FIFO[46][9] , \FIFO[46][8] ,
         \FIFO[46][7] , \FIFO[46][6] , \FIFO[46][5] , \FIFO[46][4] ,
         \FIFO[46][3] , \FIFO[46][2] , \FIFO[46][1] , \FIFO[46][0] ,
         \FIFO[47][31] , \FIFO[47][30] , \FIFO[47][29] , \FIFO[47][28] ,
         \FIFO[47][27] , \FIFO[47][26] , \FIFO[47][25] , \FIFO[47][24] ,
         \FIFO[47][23] , \FIFO[47][22] , \FIFO[47][21] , \FIFO[47][20] ,
         \FIFO[47][19] , \FIFO[47][18] , \FIFO[47][17] , \FIFO[47][16] ,
         \FIFO[47][15] , \FIFO[47][14] , \FIFO[47][13] , \FIFO[47][12] ,
         \FIFO[47][11] , \FIFO[47][10] , \FIFO[47][9] , \FIFO[47][8] ,
         \FIFO[47][7] , \FIFO[47][6] , \FIFO[47][5] , \FIFO[47][4] ,
         \FIFO[47][3] , \FIFO[47][2] , \FIFO[47][1] , \FIFO[47][0] ,
         \FIFO[48][31] , \FIFO[48][30] , \FIFO[48][29] , \FIFO[48][28] ,
         \FIFO[48][27] , \FIFO[48][26] , \FIFO[48][25] , \FIFO[48][24] ,
         \FIFO[48][23] , \FIFO[48][22] , \FIFO[48][21] , \FIFO[48][20] ,
         \FIFO[48][19] , \FIFO[48][18] , \FIFO[48][17] , \FIFO[48][16] ,
         \FIFO[48][15] , \FIFO[48][14] , \FIFO[48][13] , \FIFO[48][12] ,
         \FIFO[48][11] , \FIFO[48][10] , \FIFO[48][9] , \FIFO[48][8] ,
         \FIFO[48][7] , \FIFO[48][6] , \FIFO[48][5] , \FIFO[48][4] ,
         \FIFO[48][3] , \FIFO[48][2] , \FIFO[48][1] , \FIFO[48][0] ,
         \FIFO[49][31] , \FIFO[49][30] , \FIFO[49][29] , \FIFO[49][28] ,
         \FIFO[49][27] , \FIFO[49][26] , \FIFO[49][25] , \FIFO[49][24] ,
         \FIFO[49][23] , \FIFO[49][22] , \FIFO[49][21] , \FIFO[49][20] ,
         \FIFO[49][19] , \FIFO[49][18] , \FIFO[49][17] , \FIFO[49][16] ,
         \FIFO[49][15] , \FIFO[49][14] , \FIFO[49][13] , \FIFO[49][12] ,
         \FIFO[49][11] , \FIFO[49][10] , \FIFO[49][9] , \FIFO[49][8] ,
         \FIFO[49][7] , \FIFO[49][6] , \FIFO[49][5] , \FIFO[49][4] ,
         \FIFO[49][3] , \FIFO[49][2] , \FIFO[49][1] , \FIFO[49][0] ,
         \FIFO[50][31] , \FIFO[50][30] , \FIFO[50][29] , \FIFO[50][28] ,
         \FIFO[50][27] , \FIFO[50][26] , \FIFO[50][25] , \FIFO[50][24] ,
         \FIFO[50][23] , \FIFO[50][22] , \FIFO[50][21] , \FIFO[50][20] ,
         \FIFO[50][19] , \FIFO[50][18] , \FIFO[50][17] , \FIFO[50][16] ,
         \FIFO[50][15] , \FIFO[50][14] , \FIFO[50][13] , \FIFO[50][12] ,
         \FIFO[50][11] , \FIFO[50][10] , \FIFO[50][9] , \FIFO[50][8] ,
         \FIFO[50][7] , \FIFO[50][6] , \FIFO[50][5] , \FIFO[50][4] ,
         \FIFO[50][3] , \FIFO[50][2] , \FIFO[50][1] , \FIFO[50][0] ,
         \FIFO[51][31] , \FIFO[51][30] , \FIFO[51][29] , \FIFO[51][28] ,
         \FIFO[51][27] , \FIFO[51][26] , \FIFO[51][25] , \FIFO[51][24] ,
         \FIFO[51][23] , \FIFO[51][22] , \FIFO[51][21] , \FIFO[51][20] ,
         \FIFO[51][19] , \FIFO[51][18] , \FIFO[51][17] , \FIFO[51][16] ,
         \FIFO[51][15] , \FIFO[51][14] , \FIFO[51][13] , \FIFO[51][12] ,
         \FIFO[51][11] , \FIFO[51][10] , \FIFO[51][9] , \FIFO[51][8] ,
         \FIFO[51][7] , \FIFO[51][6] , \FIFO[51][5] , \FIFO[51][4] ,
         \FIFO[51][3] , \FIFO[51][2] , \FIFO[51][1] , \FIFO[51][0] ,
         \FIFO[52][31] , \FIFO[52][30] , \FIFO[52][29] , \FIFO[52][28] ,
         \FIFO[52][27] , \FIFO[52][26] , \FIFO[52][25] , \FIFO[52][24] ,
         \FIFO[52][23] , \FIFO[52][22] , \FIFO[52][21] , \FIFO[52][20] ,
         \FIFO[52][19] , \FIFO[52][18] , \FIFO[52][17] , \FIFO[52][16] ,
         \FIFO[52][15] , \FIFO[52][14] , \FIFO[52][13] , \FIFO[52][12] ,
         \FIFO[52][11] , \FIFO[52][10] , \FIFO[52][9] , \FIFO[52][8] ,
         \FIFO[52][7] , \FIFO[52][6] , \FIFO[52][5] , \FIFO[52][4] ,
         \FIFO[52][3] , \FIFO[52][2] , \FIFO[52][1] , \FIFO[52][0] ,
         \FIFO[53][31] , \FIFO[53][30] , \FIFO[53][29] , \FIFO[53][28] ,
         \FIFO[53][27] , \FIFO[53][26] , \FIFO[53][25] , \FIFO[53][24] ,
         \FIFO[53][23] , \FIFO[53][22] , \FIFO[53][21] , \FIFO[53][20] ,
         \FIFO[53][19] , \FIFO[53][18] , \FIFO[53][17] , \FIFO[53][16] ,
         \FIFO[53][15] , \FIFO[53][14] , \FIFO[53][13] , \FIFO[53][12] ,
         \FIFO[53][11] , \FIFO[53][10] , \FIFO[53][9] , \FIFO[53][8] ,
         \FIFO[53][7] , \FIFO[53][6] , \FIFO[53][5] , \FIFO[53][4] ,
         \FIFO[53][3] , \FIFO[53][2] , \FIFO[53][1] , \FIFO[53][0] ,
         \FIFO[54][31] , \FIFO[54][30] , \FIFO[54][29] , \FIFO[54][28] ,
         \FIFO[54][27] , \FIFO[54][26] , \FIFO[54][25] , \FIFO[54][24] ,
         \FIFO[54][23] , \FIFO[54][22] , \FIFO[54][21] , \FIFO[54][20] ,
         \FIFO[54][19] , \FIFO[54][18] , \FIFO[54][17] , \FIFO[54][16] ,
         \FIFO[54][15] , \FIFO[54][14] , \FIFO[54][13] , \FIFO[54][12] ,
         \FIFO[54][11] , \FIFO[54][10] , \FIFO[54][9] , \FIFO[54][8] ,
         \FIFO[54][7] , \FIFO[54][6] , \FIFO[54][5] , \FIFO[54][4] ,
         \FIFO[54][3] , \FIFO[54][2] , \FIFO[54][1] , \FIFO[54][0] ,
         \FIFO[55][31] , \FIFO[55][30] , \FIFO[55][29] , \FIFO[55][28] ,
         \FIFO[55][27] , \FIFO[55][26] , \FIFO[55][25] , \FIFO[55][24] ,
         \FIFO[55][23] , \FIFO[55][22] , \FIFO[55][21] , \FIFO[55][20] ,
         \FIFO[55][19] , \FIFO[55][18] , \FIFO[55][17] , \FIFO[55][16] ,
         \FIFO[55][15] , \FIFO[55][14] , \FIFO[55][13] , \FIFO[55][12] ,
         \FIFO[55][11] , \FIFO[55][10] , \FIFO[55][9] , \FIFO[55][8] ,
         \FIFO[55][7] , \FIFO[55][6] , \FIFO[55][5] , \FIFO[55][4] ,
         \FIFO[55][3] , \FIFO[55][2] , \FIFO[55][1] , \FIFO[55][0] ,
         \FIFO[56][31] , \FIFO[56][30] , \FIFO[56][29] , \FIFO[56][28] ,
         \FIFO[56][27] , \FIFO[56][26] , \FIFO[56][25] , \FIFO[56][24] ,
         \FIFO[56][23] , \FIFO[56][22] , \FIFO[56][21] , \FIFO[56][20] ,
         \FIFO[56][19] , \FIFO[56][18] , \FIFO[56][17] , \FIFO[56][16] ,
         \FIFO[56][15] , \FIFO[56][14] , \FIFO[56][13] , \FIFO[56][12] ,
         \FIFO[56][11] , \FIFO[56][10] , \FIFO[56][9] , \FIFO[56][8] ,
         \FIFO[56][7] , \FIFO[56][6] , \FIFO[56][5] , \FIFO[56][4] ,
         \FIFO[56][3] , \FIFO[56][2] , \FIFO[56][1] , \FIFO[56][0] ,
         \FIFO[57][31] , \FIFO[57][30] , \FIFO[57][29] , \FIFO[57][28] ,
         \FIFO[57][27] , \FIFO[57][26] , \FIFO[57][25] , \FIFO[57][24] ,
         \FIFO[57][23] , \FIFO[57][22] , \FIFO[57][21] , \FIFO[57][20] ,
         \FIFO[57][19] , \FIFO[57][18] , \FIFO[57][17] , \FIFO[57][16] ,
         \FIFO[57][15] , \FIFO[57][14] , \FIFO[57][13] , \FIFO[57][12] ,
         \FIFO[57][11] , \FIFO[57][10] , \FIFO[57][9] , \FIFO[57][8] ,
         \FIFO[57][7] , \FIFO[57][6] , \FIFO[57][5] , \FIFO[57][4] ,
         \FIFO[57][3] , \FIFO[57][2] , \FIFO[57][1] , \FIFO[57][0] ,
         \FIFO[58][31] , \FIFO[58][30] , \FIFO[58][29] , \FIFO[58][28] ,
         \FIFO[58][27] , \FIFO[58][26] , \FIFO[58][25] , \FIFO[58][24] ,
         \FIFO[58][23] , \FIFO[58][22] , \FIFO[58][21] , \FIFO[58][20] ,
         \FIFO[58][19] , \FIFO[58][18] , \FIFO[58][17] , \FIFO[58][16] ,
         \FIFO[58][15] , \FIFO[58][14] , \FIFO[58][13] , \FIFO[58][12] ,
         \FIFO[58][11] , \FIFO[58][10] , \FIFO[58][9] , \FIFO[58][8] ,
         \FIFO[58][7] , \FIFO[58][6] , \FIFO[58][5] , \FIFO[58][4] ,
         \FIFO[58][3] , \FIFO[58][2] , \FIFO[58][1] , \FIFO[58][0] ,
         \FIFO[59][31] , \FIFO[59][30] , \FIFO[59][29] , \FIFO[59][28] ,
         \FIFO[59][27] , \FIFO[59][26] , \FIFO[59][25] , \FIFO[59][24] ,
         \FIFO[59][23] , \FIFO[59][22] , \FIFO[59][21] , \FIFO[59][20] ,
         \FIFO[59][19] , \FIFO[59][18] , \FIFO[59][17] , \FIFO[59][16] ,
         \FIFO[59][15] , \FIFO[59][14] , \FIFO[59][13] , \FIFO[59][12] ,
         \FIFO[59][11] , \FIFO[59][10] , \FIFO[59][9] , \FIFO[59][8] ,
         \FIFO[59][7] , \FIFO[59][6] , \FIFO[59][5] , \FIFO[59][4] ,
         \FIFO[59][3] , \FIFO[59][2] , \FIFO[59][1] , \FIFO[59][0] ,
         \FIFO[60][31] , \FIFO[60][30] , \FIFO[60][29] , \FIFO[60][28] ,
         \FIFO[60][27] , \FIFO[60][26] , \FIFO[60][25] , \FIFO[60][24] ,
         \FIFO[60][23] , \FIFO[60][22] , \FIFO[60][21] , \FIFO[60][20] ,
         \FIFO[60][19] , \FIFO[60][18] , \FIFO[60][17] , \FIFO[60][16] ,
         \FIFO[60][15] , \FIFO[60][14] , \FIFO[60][13] , \FIFO[60][12] ,
         \FIFO[60][11] , \FIFO[60][10] , \FIFO[60][9] , \FIFO[60][8] ,
         \FIFO[60][7] , \FIFO[60][6] , \FIFO[60][5] , \FIFO[60][4] ,
         \FIFO[60][3] , \FIFO[60][2] , \FIFO[60][1] , \FIFO[60][0] ,
         \FIFO[61][31] , \FIFO[61][30] , \FIFO[61][29] , \FIFO[61][28] ,
         \FIFO[61][27] , \FIFO[61][26] , \FIFO[61][25] , \FIFO[61][24] ,
         \FIFO[61][23] , \FIFO[61][22] , \FIFO[61][21] , \FIFO[61][20] ,
         \FIFO[61][19] , \FIFO[61][18] , \FIFO[61][17] , \FIFO[61][16] ,
         \FIFO[61][15] , \FIFO[61][14] , \FIFO[61][13] , \FIFO[61][12] ,
         \FIFO[61][11] , \FIFO[61][10] , \FIFO[61][9] , \FIFO[61][8] ,
         \FIFO[61][7] , \FIFO[61][6] , \FIFO[61][5] , \FIFO[61][4] ,
         \FIFO[61][3] , \FIFO[61][2] , \FIFO[61][1] , \FIFO[61][0] ,
         \FIFO[62][31] , \FIFO[62][30] , \FIFO[62][29] , \FIFO[62][28] ,
         \FIFO[62][27] , \FIFO[62][26] , \FIFO[62][25] , \FIFO[62][24] ,
         \FIFO[62][23] , \FIFO[62][22] , \FIFO[62][21] , \FIFO[62][20] ,
         \FIFO[62][19] , \FIFO[62][18] , \FIFO[62][17] , \FIFO[62][16] ,
         \FIFO[62][15] , \FIFO[62][14] , \FIFO[62][13] , \FIFO[62][12] ,
         \FIFO[62][11] , \FIFO[62][10] , \FIFO[62][9] , \FIFO[62][8] ,
         \FIFO[62][7] , \FIFO[62][6] , \FIFO[62][5] , \FIFO[62][4] ,
         \FIFO[62][3] , \FIFO[62][2] , \FIFO[62][1] , \FIFO[62][0] ,
         \FIFO[63][31] , \FIFO[63][30] , \FIFO[63][29] , \FIFO[63][28] ,
         \FIFO[63][27] , \FIFO[63][26] , \FIFO[63][25] , \FIFO[63][24] ,
         \FIFO[63][23] , \FIFO[63][22] , \FIFO[63][21] , \FIFO[63][20] ,
         \FIFO[63][19] , \FIFO[63][18] , \FIFO[63][17] , \FIFO[63][16] ,
         \FIFO[63][15] , \FIFO[63][14] , \FIFO[63][13] , \FIFO[63][12] ,
         \FIFO[63][11] , \FIFO[63][10] , \FIFO[63][9] , \FIFO[63][8] ,
         \FIFO[63][7] , \FIFO[63][6] , \FIFO[63][5] , \FIFO[63][4] ,
         \FIFO[63][3] , \FIFO[63][2] , \FIFO[63][1] , \FIFO[63][0] ,
         \FIFO[64][31] , \FIFO[64][30] , \FIFO[64][29] , \FIFO[64][28] ,
         \FIFO[64][27] , \FIFO[64][26] , \FIFO[64][25] , \FIFO[64][24] ,
         \FIFO[64][23] , \FIFO[64][22] , \FIFO[64][21] , \FIFO[64][20] ,
         \FIFO[64][19] , \FIFO[64][18] , \FIFO[64][17] , \FIFO[64][16] ,
         \FIFO[64][15] , \FIFO[64][14] , \FIFO[64][13] , \FIFO[64][12] ,
         \FIFO[64][11] , \FIFO[64][10] , \FIFO[64][9] , \FIFO[64][8] ,
         \FIFO[64][7] , \FIFO[64][6] , \FIFO[64][5] , \FIFO[64][4] ,
         \FIFO[64][3] , \FIFO[64][2] , \FIFO[64][1] , \FIFO[64][0] ,
         \FIFO[65][31] , \FIFO[65][30] , \FIFO[65][29] , \FIFO[65][28] ,
         \FIFO[65][27] , \FIFO[65][26] , \FIFO[65][25] , \FIFO[65][24] ,
         \FIFO[65][23] , \FIFO[65][22] , \FIFO[65][21] , \FIFO[65][20] ,
         \FIFO[65][19] , \FIFO[65][18] , \FIFO[65][17] , \FIFO[65][16] ,
         \FIFO[65][15] , \FIFO[65][14] , \FIFO[65][13] , \FIFO[65][12] ,
         \FIFO[65][11] , \FIFO[65][10] , \FIFO[65][9] , \FIFO[65][8] ,
         \FIFO[65][7] , \FIFO[65][6] , \FIFO[65][5] , \FIFO[65][4] ,
         \FIFO[65][3] , \FIFO[65][2] , \FIFO[65][1] , \FIFO[65][0] ,
         \FIFO[66][31] , \FIFO[66][30] , \FIFO[66][29] , \FIFO[66][28] ,
         \FIFO[66][27] , \FIFO[66][26] , \FIFO[66][25] , \FIFO[66][24] ,
         \FIFO[66][23] , \FIFO[66][22] , \FIFO[66][21] , \FIFO[66][20] ,
         \FIFO[66][19] , \FIFO[66][18] , \FIFO[66][17] , \FIFO[66][16] ,
         \FIFO[66][15] , \FIFO[66][14] , \FIFO[66][13] , \FIFO[66][12] ,
         \FIFO[66][11] , \FIFO[66][10] , \FIFO[66][9] , \FIFO[66][8] ,
         \FIFO[66][7] , \FIFO[66][6] , \FIFO[66][5] , \FIFO[66][4] ,
         \FIFO[66][3] , \FIFO[66][2] , \FIFO[66][1] , \FIFO[66][0] ,
         \FIFO[67][31] , \FIFO[67][30] , \FIFO[67][29] , \FIFO[67][28] ,
         \FIFO[67][27] , \FIFO[67][26] , \FIFO[67][25] , \FIFO[67][24] ,
         \FIFO[67][23] , \FIFO[67][22] , \FIFO[67][21] , \FIFO[67][20] ,
         \FIFO[67][19] , \FIFO[67][18] , \FIFO[67][17] , \FIFO[67][16] ,
         \FIFO[67][15] , \FIFO[67][14] , \FIFO[67][13] , \FIFO[67][12] ,
         \FIFO[67][11] , \FIFO[67][10] , \FIFO[67][9] , \FIFO[67][8] ,
         \FIFO[67][7] , \FIFO[67][6] , \FIFO[67][5] , \FIFO[67][4] ,
         \FIFO[67][3] , \FIFO[67][2] , \FIFO[67][1] , \FIFO[67][0] ,
         \FIFO[68][31] , \FIFO[68][30] , \FIFO[68][29] , \FIFO[68][28] ,
         \FIFO[68][27] , \FIFO[68][26] , \FIFO[68][25] , \FIFO[68][24] ,
         \FIFO[68][23] , \FIFO[68][22] , \FIFO[68][21] , \FIFO[68][20] ,
         \FIFO[68][19] , \FIFO[68][18] , \FIFO[68][17] , \FIFO[68][16] ,
         \FIFO[68][15] , \FIFO[68][14] , \FIFO[68][13] , \FIFO[68][12] ,
         \FIFO[68][11] , \FIFO[68][10] , \FIFO[68][9] , \FIFO[68][8] ,
         \FIFO[68][7] , \FIFO[68][6] , \FIFO[68][5] , \FIFO[68][4] ,
         \FIFO[68][3] , \FIFO[68][2] , \FIFO[68][1] , \FIFO[68][0] ,
         \FIFO[69][31] , \FIFO[69][30] , \FIFO[69][29] , \FIFO[69][28] ,
         \FIFO[69][27] , \FIFO[69][26] , \FIFO[69][25] , \FIFO[69][24] ,
         \FIFO[69][23] , \FIFO[69][22] , \FIFO[69][21] , \FIFO[69][20] ,
         \FIFO[69][19] , \FIFO[69][18] , \FIFO[69][17] , \FIFO[69][16] ,
         \FIFO[69][15] , \FIFO[69][14] , \FIFO[69][13] , \FIFO[69][12] ,
         \FIFO[69][11] , \FIFO[69][10] , \FIFO[69][9] , \FIFO[69][8] ,
         \FIFO[69][7] , \FIFO[69][6] , \FIFO[69][5] , \FIFO[69][4] ,
         \FIFO[69][3] , \FIFO[69][2] , \FIFO[69][1] , \FIFO[69][0] ,
         \FIFO[70][31] , \FIFO[70][30] , \FIFO[70][29] , \FIFO[70][28] ,
         \FIFO[70][27] , \FIFO[70][26] , \FIFO[70][25] , \FIFO[70][24] ,
         \FIFO[70][23] , \FIFO[70][22] , \FIFO[70][21] , \FIFO[70][20] ,
         \FIFO[70][19] , \FIFO[70][18] , \FIFO[70][17] , \FIFO[70][16] ,
         \FIFO[70][15] , \FIFO[70][14] , \FIFO[70][13] , \FIFO[70][12] ,
         \FIFO[70][11] , \FIFO[70][10] , \FIFO[70][9] , \FIFO[70][8] ,
         \FIFO[70][7] , \FIFO[70][6] , \FIFO[70][5] , \FIFO[70][4] ,
         \FIFO[70][3] , \FIFO[70][2] , \FIFO[70][1] , \FIFO[70][0] ,
         \FIFO[71][31] , \FIFO[71][30] , \FIFO[71][29] , \FIFO[71][28] ,
         \FIFO[71][27] , \FIFO[71][26] , \FIFO[71][25] , \FIFO[71][24] ,
         \FIFO[71][23] , \FIFO[71][22] , \FIFO[71][21] , \FIFO[71][20] ,
         \FIFO[71][19] , \FIFO[71][18] , \FIFO[71][17] , \FIFO[71][16] ,
         \FIFO[71][15] , \FIFO[71][14] , \FIFO[71][13] , \FIFO[71][12] ,
         \FIFO[71][11] , \FIFO[71][10] , \FIFO[71][9] , \FIFO[71][8] ,
         \FIFO[71][7] , \FIFO[71][6] , \FIFO[71][5] , \FIFO[71][4] ,
         \FIFO[71][3] , \FIFO[71][2] , \FIFO[71][1] , \FIFO[71][0] ,
         \FIFO[72][31] , \FIFO[72][30] , \FIFO[72][29] , \FIFO[72][28] ,
         \FIFO[72][27] , \FIFO[72][26] , \FIFO[72][25] , \FIFO[72][24] ,
         \FIFO[72][23] , \FIFO[72][22] , \FIFO[72][21] , \FIFO[72][20] ,
         \FIFO[72][19] , \FIFO[72][18] , \FIFO[72][17] , \FIFO[72][16] ,
         \FIFO[72][15] , \FIFO[72][14] , \FIFO[72][13] , \FIFO[72][12] ,
         \FIFO[72][11] , \FIFO[72][10] , \FIFO[72][9] , \FIFO[72][8] ,
         \FIFO[72][7] , \FIFO[72][6] , \FIFO[72][5] , \FIFO[72][4] ,
         \FIFO[72][3] , \FIFO[72][2] , \FIFO[72][1] , \FIFO[72][0] ,
         \FIFO[73][31] , \FIFO[73][30] , \FIFO[73][29] , \FIFO[73][28] ,
         \FIFO[73][27] , \FIFO[73][26] , \FIFO[73][25] , \FIFO[73][24] ,
         \FIFO[73][23] , \FIFO[73][22] , \FIFO[73][21] , \FIFO[73][20] ,
         \FIFO[73][19] , \FIFO[73][18] , \FIFO[73][17] , \FIFO[73][16] ,
         \FIFO[73][15] , \FIFO[73][14] , \FIFO[73][13] , \FIFO[73][12] ,
         \FIFO[73][11] , \FIFO[73][10] , \FIFO[73][9] , \FIFO[73][8] ,
         \FIFO[73][7] , \FIFO[73][6] , \FIFO[73][5] , \FIFO[73][4] ,
         \FIFO[73][3] , \FIFO[73][2] , \FIFO[73][1] , \FIFO[73][0] ,
         \FIFO[74][31] , \FIFO[74][30] , \FIFO[74][29] , \FIFO[74][28] ,
         \FIFO[74][27] , \FIFO[74][26] , \FIFO[74][25] , \FIFO[74][24] ,
         \FIFO[74][23] , \FIFO[74][22] , \FIFO[74][21] , \FIFO[74][20] ,
         \FIFO[74][19] , \FIFO[74][18] , \FIFO[74][17] , \FIFO[74][16] ,
         \FIFO[74][15] , \FIFO[74][14] , \FIFO[74][13] , \FIFO[74][12] ,
         \FIFO[74][11] , \FIFO[74][10] , \FIFO[74][9] , \FIFO[74][8] ,
         \FIFO[74][7] , \FIFO[74][6] , \FIFO[74][5] , \FIFO[74][4] ,
         \FIFO[74][3] , \FIFO[74][2] , \FIFO[74][1] , \FIFO[74][0] ,
         \FIFO[75][31] , \FIFO[75][30] , \FIFO[75][29] , \FIFO[75][28] ,
         \FIFO[75][27] , \FIFO[75][26] , \FIFO[75][25] , \FIFO[75][24] ,
         \FIFO[75][23] , \FIFO[75][22] , \FIFO[75][21] , \FIFO[75][20] ,
         \FIFO[75][19] , \FIFO[75][18] , \FIFO[75][17] , \FIFO[75][16] ,
         \FIFO[75][15] , \FIFO[75][14] , \FIFO[75][13] , \FIFO[75][12] ,
         \FIFO[75][11] , \FIFO[75][10] , \FIFO[75][9] , \FIFO[75][8] ,
         \FIFO[75][7] , \FIFO[75][6] , \FIFO[75][5] , \FIFO[75][4] ,
         \FIFO[75][3] , \FIFO[75][2] , \FIFO[75][1] , \FIFO[75][0] ,
         \FIFO[76][31] , \FIFO[76][30] , \FIFO[76][29] , \FIFO[76][28] ,
         \FIFO[76][27] , \FIFO[76][26] , \FIFO[76][25] , \FIFO[76][24] ,
         \FIFO[76][23] , \FIFO[76][22] , \FIFO[76][21] , \FIFO[76][20] ,
         \FIFO[76][19] , \FIFO[76][18] , \FIFO[76][17] , \FIFO[76][16] ,
         \FIFO[76][15] , \FIFO[76][14] , \FIFO[76][13] , \FIFO[76][12] ,
         \FIFO[76][11] , \FIFO[76][10] , \FIFO[76][9] , \FIFO[76][8] ,
         \FIFO[76][7] , \FIFO[76][6] , \FIFO[76][5] , \FIFO[76][4] ,
         \FIFO[76][3] , \FIFO[76][2] , \FIFO[76][1] , \FIFO[76][0] ,
         \FIFO[77][31] , \FIFO[77][30] , \FIFO[77][29] , \FIFO[77][28] ,
         \FIFO[77][27] , \FIFO[77][26] , \FIFO[77][25] , \FIFO[77][24] ,
         \FIFO[77][23] , \FIFO[77][22] , \FIFO[77][21] , \FIFO[77][20] ,
         \FIFO[77][19] , \FIFO[77][18] , \FIFO[77][17] , \FIFO[77][16] ,
         \FIFO[77][15] , \FIFO[77][14] , \FIFO[77][13] , \FIFO[77][12] ,
         \FIFO[77][11] , \FIFO[77][10] , \FIFO[77][9] , \FIFO[77][8] ,
         \FIFO[77][7] , \FIFO[77][6] , \FIFO[77][5] , \FIFO[77][4] ,
         \FIFO[77][3] , \FIFO[77][2] , \FIFO[77][1] , \FIFO[77][0] ,
         \FIFO[78][31] , \FIFO[78][30] , \FIFO[78][29] , \FIFO[78][28] ,
         \FIFO[78][27] , \FIFO[78][26] , \FIFO[78][25] , \FIFO[78][24] ,
         \FIFO[78][23] , \FIFO[78][22] , \FIFO[78][21] , \FIFO[78][20] ,
         \FIFO[78][19] , \FIFO[78][18] , \FIFO[78][17] , \FIFO[78][16] ,
         \FIFO[78][15] , \FIFO[78][14] , \FIFO[78][13] , \FIFO[78][12] ,
         \FIFO[78][11] , \FIFO[78][10] , \FIFO[78][9] , \FIFO[78][8] ,
         \FIFO[78][7] , \FIFO[78][6] , \FIFO[78][5] , \FIFO[78][4] ,
         \FIFO[78][3] , \FIFO[78][2] , \FIFO[78][1] , \FIFO[78][0] ,
         \FIFO[79][31] , \FIFO[79][30] , \FIFO[79][29] , \FIFO[79][28] ,
         \FIFO[79][27] , \FIFO[79][26] , \FIFO[79][25] , \FIFO[79][24] ,
         \FIFO[79][23] , \FIFO[79][22] , \FIFO[79][21] , \FIFO[79][20] ,
         \FIFO[79][19] , \FIFO[79][18] , \FIFO[79][17] , \FIFO[79][16] ,
         \FIFO[79][15] , \FIFO[79][14] , \FIFO[79][13] , \FIFO[79][12] ,
         \FIFO[79][11] , \FIFO[79][10] , \FIFO[79][9] , \FIFO[79][8] ,
         \FIFO[79][7] , \FIFO[79][6] , \FIFO[79][5] , \FIFO[79][4] ,
         \FIFO[79][3] , \FIFO[79][2] , \FIFO[79][1] , \FIFO[79][0] ,
         \FIFO[80][31] , \FIFO[80][30] , \FIFO[80][29] , \FIFO[80][28] ,
         \FIFO[80][27] , \FIFO[80][26] , \FIFO[80][25] , \FIFO[80][24] ,
         \FIFO[80][23] , \FIFO[80][22] , \FIFO[80][21] , \FIFO[80][20] ,
         \FIFO[80][19] , \FIFO[80][18] , \FIFO[80][17] , \FIFO[80][16] ,
         \FIFO[80][15] , \FIFO[80][14] , \FIFO[80][13] , \FIFO[80][12] ,
         \FIFO[80][11] , \FIFO[80][10] , \FIFO[80][9] , \FIFO[80][8] ,
         \FIFO[80][7] , \FIFO[80][6] , \FIFO[80][5] , \FIFO[80][4] ,
         \FIFO[80][3] , \FIFO[80][2] , \FIFO[80][1] , \FIFO[80][0] ,
         \FIFO[81][31] , \FIFO[81][30] , \FIFO[81][29] , \FIFO[81][28] ,
         \FIFO[81][27] , \FIFO[81][26] , \FIFO[81][25] , \FIFO[81][24] ,
         \FIFO[81][23] , \FIFO[81][22] , \FIFO[81][21] , \FIFO[81][20] ,
         \FIFO[81][19] , \FIFO[81][18] , \FIFO[81][17] , \FIFO[81][16] ,
         \FIFO[81][15] , \FIFO[81][14] , \FIFO[81][13] , \FIFO[81][12] ,
         \FIFO[81][11] , \FIFO[81][10] , \FIFO[81][9] , \FIFO[81][8] ,
         \FIFO[81][7] , \FIFO[81][6] , \FIFO[81][5] , \FIFO[81][4] ,
         \FIFO[81][3] , \FIFO[81][2] , \FIFO[81][1] , \FIFO[81][0] ,
         \FIFO[82][31] , \FIFO[82][30] , \FIFO[82][29] , \FIFO[82][28] ,
         \FIFO[82][27] , \FIFO[82][26] , \FIFO[82][25] , \FIFO[82][24] ,
         \FIFO[82][23] , \FIFO[82][22] , \FIFO[82][21] , \FIFO[82][20] ,
         \FIFO[82][19] , \FIFO[82][18] , \FIFO[82][17] , \FIFO[82][16] ,
         \FIFO[82][15] , \FIFO[82][14] , \FIFO[82][13] , \FIFO[82][12] ,
         \FIFO[82][11] , \FIFO[82][10] , \FIFO[82][9] , \FIFO[82][8] ,
         \FIFO[82][7] , \FIFO[82][6] , \FIFO[82][5] , \FIFO[82][4] ,
         \FIFO[82][3] , \FIFO[82][2] , \FIFO[82][1] , \FIFO[82][0] ,
         \FIFO[83][31] , \FIFO[83][30] , \FIFO[83][29] , \FIFO[83][28] ,
         \FIFO[83][27] , \FIFO[83][26] , \FIFO[83][25] , \FIFO[83][24] ,
         \FIFO[83][23] , \FIFO[83][22] , \FIFO[83][21] , \FIFO[83][20] ,
         \FIFO[83][19] , \FIFO[83][18] , \FIFO[83][17] , \FIFO[83][16] ,
         \FIFO[83][15] , \FIFO[83][14] , \FIFO[83][13] , \FIFO[83][12] ,
         \FIFO[83][11] , \FIFO[83][10] , \FIFO[83][9] , \FIFO[83][8] ,
         \FIFO[83][7] , \FIFO[83][6] , \FIFO[83][5] , \FIFO[83][4] ,
         \FIFO[83][3] , \FIFO[83][2] , \FIFO[83][1] , \FIFO[83][0] ,
         \FIFO[84][31] , \FIFO[84][30] , \FIFO[84][29] , \FIFO[84][28] ,
         \FIFO[84][27] , \FIFO[84][26] , \FIFO[84][25] , \FIFO[84][24] ,
         \FIFO[84][23] , \FIFO[84][22] , \FIFO[84][21] , \FIFO[84][20] ,
         \FIFO[84][19] , \FIFO[84][18] , \FIFO[84][17] , \FIFO[84][16] ,
         \FIFO[84][15] , \FIFO[84][14] , \FIFO[84][13] , \FIFO[84][12] ,
         \FIFO[84][11] , \FIFO[84][10] , \FIFO[84][9] , \FIFO[84][8] ,
         \FIFO[84][7] , \FIFO[84][6] , \FIFO[84][5] , \FIFO[84][4] ,
         \FIFO[84][3] , \FIFO[84][2] , \FIFO[84][1] , \FIFO[84][0] ,
         \FIFO[85][31] , \FIFO[85][30] , \FIFO[85][29] , \FIFO[85][28] ,
         \FIFO[85][27] , \FIFO[85][26] , \FIFO[85][25] , \FIFO[85][24] ,
         \FIFO[85][23] , \FIFO[85][22] , \FIFO[85][21] , \FIFO[85][20] ,
         \FIFO[85][19] , \FIFO[85][18] , \FIFO[85][17] , \FIFO[85][16] ,
         \FIFO[85][15] , \FIFO[85][14] , \FIFO[85][13] , \FIFO[85][12] ,
         \FIFO[85][11] , \FIFO[85][10] , \FIFO[85][9] , \FIFO[85][8] ,
         \FIFO[85][7] , \FIFO[85][6] , \FIFO[85][5] , \FIFO[85][4] ,
         \FIFO[85][3] , \FIFO[85][2] , \FIFO[85][1] , \FIFO[85][0] ,
         \FIFO[86][31] , \FIFO[86][30] , \FIFO[86][29] , \FIFO[86][28] ,
         \FIFO[86][27] , \FIFO[86][26] , \FIFO[86][25] , \FIFO[86][24] ,
         \FIFO[86][23] , \FIFO[86][22] , \FIFO[86][21] , \FIFO[86][20] ,
         \FIFO[86][19] , \FIFO[86][18] , \FIFO[86][17] , \FIFO[86][16] ,
         \FIFO[86][15] , \FIFO[86][14] , \FIFO[86][13] , \FIFO[86][12] ,
         \FIFO[86][11] , \FIFO[86][10] , \FIFO[86][9] , \FIFO[86][8] ,
         \FIFO[86][7] , \FIFO[86][6] , \FIFO[86][5] , \FIFO[86][4] ,
         \FIFO[86][3] , \FIFO[86][2] , \FIFO[86][1] , \FIFO[86][0] ,
         \FIFO[87][31] , \FIFO[87][30] , \FIFO[87][29] , \FIFO[87][28] ,
         \FIFO[87][27] , \FIFO[87][26] , \FIFO[87][25] , \FIFO[87][24] ,
         \FIFO[87][23] , \FIFO[87][22] , \FIFO[87][21] , \FIFO[87][20] ,
         \FIFO[87][19] , \FIFO[87][18] , \FIFO[87][17] , \FIFO[87][16] ,
         \FIFO[87][15] , \FIFO[87][14] , \FIFO[87][13] , \FIFO[87][12] ,
         \FIFO[87][11] , \FIFO[87][10] , \FIFO[87][9] , \FIFO[87][8] ,
         \FIFO[87][7] , \FIFO[87][6] , \FIFO[87][5] , \FIFO[87][4] ,
         \FIFO[87][3] , \FIFO[87][2] , \FIFO[87][1] , \FIFO[87][0] ,
         \FIFO[88][31] , \FIFO[88][30] , \FIFO[88][29] , \FIFO[88][28] ,
         \FIFO[88][27] , \FIFO[88][26] , \FIFO[88][25] , \FIFO[88][24] ,
         \FIFO[88][23] , \FIFO[88][22] , \FIFO[88][21] , \FIFO[88][20] ,
         \FIFO[88][19] , \FIFO[88][18] , \FIFO[88][17] , \FIFO[88][16] ,
         \FIFO[88][15] , \FIFO[88][14] , \FIFO[88][13] , \FIFO[88][12] ,
         \FIFO[88][11] , \FIFO[88][10] , \FIFO[88][9] , \FIFO[88][8] ,
         \FIFO[88][7] , \FIFO[88][6] , \FIFO[88][5] , \FIFO[88][4] ,
         \FIFO[88][3] , \FIFO[88][2] , \FIFO[88][1] , \FIFO[88][0] ,
         \FIFO[89][31] , \FIFO[89][30] , \FIFO[89][29] , \FIFO[89][28] ,
         \FIFO[89][27] , \FIFO[89][26] , \FIFO[89][25] , \FIFO[89][24] ,
         \FIFO[89][23] , \FIFO[89][22] , \FIFO[89][21] , \FIFO[89][20] ,
         \FIFO[89][19] , \FIFO[89][18] , \FIFO[89][17] , \FIFO[89][16] ,
         \FIFO[89][15] , \FIFO[89][14] , \FIFO[89][13] , \FIFO[89][12] ,
         \FIFO[89][11] , \FIFO[89][10] , \FIFO[89][9] , \FIFO[89][8] ,
         \FIFO[89][7] , \FIFO[89][6] , \FIFO[89][5] , \FIFO[89][4] ,
         \FIFO[89][3] , \FIFO[89][2] , \FIFO[89][1] , \FIFO[89][0] ,
         \FIFO[90][31] , \FIFO[90][30] , \FIFO[90][29] , \FIFO[90][28] ,
         \FIFO[90][27] , \FIFO[90][26] , \FIFO[90][25] , \FIFO[90][24] ,
         \FIFO[90][23] , \FIFO[90][22] , \FIFO[90][21] , \FIFO[90][20] ,
         \FIFO[90][19] , \FIFO[90][18] , \FIFO[90][17] , \FIFO[90][16] ,
         \FIFO[90][15] , \FIFO[90][14] , \FIFO[90][13] , \FIFO[90][12] ,
         \FIFO[90][11] , \FIFO[90][10] , \FIFO[90][9] , \FIFO[90][8] ,
         \FIFO[90][7] , \FIFO[90][6] , \FIFO[90][5] , \FIFO[90][4] ,
         \FIFO[90][3] , \FIFO[90][2] , \FIFO[90][1] , \FIFO[90][0] ,
         \FIFO[91][31] , \FIFO[91][30] , \FIFO[91][29] , \FIFO[91][28] ,
         \FIFO[91][27] , \FIFO[91][26] , \FIFO[91][25] , \FIFO[91][24] ,
         \FIFO[91][23] , \FIFO[91][22] , \FIFO[91][21] , \FIFO[91][20] ,
         \FIFO[91][19] , \FIFO[91][18] , \FIFO[91][17] , \FIFO[91][16] ,
         \FIFO[91][15] , \FIFO[91][14] , \FIFO[91][13] , \FIFO[91][12] ,
         \FIFO[91][11] , \FIFO[91][10] , \FIFO[91][9] , \FIFO[91][8] ,
         \FIFO[91][7] , \FIFO[91][6] , \FIFO[91][5] , \FIFO[91][4] ,
         \FIFO[91][3] , \FIFO[91][2] , \FIFO[91][1] , \FIFO[91][0] ,
         \FIFO[92][31] , \FIFO[92][30] , \FIFO[92][29] , \FIFO[92][28] ,
         \FIFO[92][27] , \FIFO[92][26] , \FIFO[92][25] , \FIFO[92][24] ,
         \FIFO[92][23] , \FIFO[92][22] , \FIFO[92][21] , \FIFO[92][20] ,
         \FIFO[92][19] , \FIFO[92][18] , \FIFO[92][17] , \FIFO[92][16] ,
         \FIFO[92][15] , \FIFO[92][14] , \FIFO[92][13] , \FIFO[92][12] ,
         \FIFO[92][11] , \FIFO[92][10] , \FIFO[92][9] , \FIFO[92][8] ,
         \FIFO[92][7] , \FIFO[92][6] , \FIFO[92][5] , \FIFO[92][4] ,
         \FIFO[92][3] , \FIFO[92][2] , \FIFO[92][1] , \FIFO[92][0] ,
         \FIFO[93][31] , \FIFO[93][30] , \FIFO[93][29] , \FIFO[93][28] ,
         \FIFO[93][27] , \FIFO[93][26] , \FIFO[93][25] , \FIFO[93][24] ,
         \FIFO[93][23] , \FIFO[93][22] , \FIFO[93][21] , \FIFO[93][20] ,
         \FIFO[93][19] , \FIFO[93][18] , \FIFO[93][17] , \FIFO[93][16] ,
         \FIFO[93][15] , \FIFO[93][14] , \FIFO[93][13] , \FIFO[93][12] ,
         \FIFO[93][11] , \FIFO[93][10] , \FIFO[93][9] , \FIFO[93][8] ,
         \FIFO[93][7] , \FIFO[93][6] , \FIFO[93][5] , \FIFO[93][4] ,
         \FIFO[93][3] , \FIFO[93][2] , \FIFO[93][1] , \FIFO[93][0] ,
         \FIFO[94][31] , \FIFO[94][30] , \FIFO[94][29] , \FIFO[94][28] ,
         \FIFO[94][27] , \FIFO[94][26] , \FIFO[94][25] , \FIFO[94][24] ,
         \FIFO[94][23] , \FIFO[94][22] , \FIFO[94][21] , \FIFO[94][20] ,
         \FIFO[94][19] , \FIFO[94][18] , \FIFO[94][17] , \FIFO[94][16] ,
         \FIFO[94][15] , \FIFO[94][14] , \FIFO[94][13] , \FIFO[94][12] ,
         \FIFO[94][11] , \FIFO[94][10] , \FIFO[94][9] , \FIFO[94][8] ,
         \FIFO[94][7] , \FIFO[94][6] , \FIFO[94][5] , \FIFO[94][4] ,
         \FIFO[94][3] , \FIFO[94][2] , \FIFO[94][1] , \FIFO[94][0] ,
         \FIFO[95][31] , \FIFO[95][30] , \FIFO[95][29] , \FIFO[95][28] ,
         \FIFO[95][27] , \FIFO[95][26] , \FIFO[95][25] , \FIFO[95][24] ,
         \FIFO[95][23] , \FIFO[95][22] , \FIFO[95][21] , \FIFO[95][20] ,
         \FIFO[95][19] , \FIFO[95][18] , \FIFO[95][17] , \FIFO[95][16] ,
         \FIFO[95][15] , \FIFO[95][14] , \FIFO[95][13] , \FIFO[95][12] ,
         \FIFO[95][11] , \FIFO[95][10] , \FIFO[95][9] , \FIFO[95][8] ,
         \FIFO[95][7] , \FIFO[95][6] , \FIFO[95][5] , \FIFO[95][4] ,
         \FIFO[95][3] , \FIFO[95][2] , \FIFO[95][1] , \FIFO[95][0] ,
         \FIFO[96][31] , \FIFO[96][30] , \FIFO[96][29] , \FIFO[96][28] ,
         \FIFO[96][27] , \FIFO[96][26] , \FIFO[96][25] , \FIFO[96][24] ,
         \FIFO[96][23] , \FIFO[96][22] , \FIFO[96][21] , \FIFO[96][20] ,
         \FIFO[96][19] , \FIFO[96][18] , \FIFO[96][17] , \FIFO[96][16] ,
         \FIFO[96][15] , \FIFO[96][14] , \FIFO[96][13] , \FIFO[96][12] ,
         \FIFO[96][11] , \FIFO[96][10] , \FIFO[96][9] , \FIFO[96][8] ,
         \FIFO[96][7] , \FIFO[96][6] , \FIFO[96][5] , \FIFO[96][4] ,
         \FIFO[96][3] , \FIFO[96][2] , \FIFO[96][1] , \FIFO[96][0] ,
         \FIFO[97][31] , \FIFO[97][30] , \FIFO[97][29] , \FIFO[97][28] ,
         \FIFO[97][27] , \FIFO[97][26] , \FIFO[97][25] , \FIFO[97][24] ,
         \FIFO[97][23] , \FIFO[97][22] , \FIFO[97][21] , \FIFO[97][20] ,
         \FIFO[97][19] , \FIFO[97][18] , \FIFO[97][17] , \FIFO[97][16] ,
         \FIFO[97][15] , \FIFO[97][14] , \FIFO[97][13] , \FIFO[97][12] ,
         \FIFO[97][11] , \FIFO[97][10] , \FIFO[97][9] , \FIFO[97][8] ,
         \FIFO[97][7] , \FIFO[97][6] , \FIFO[97][5] , \FIFO[97][4] ,
         \FIFO[97][3] , \FIFO[97][2] , \FIFO[97][1] , \FIFO[97][0] ,
         \FIFO[98][31] , \FIFO[98][30] , \FIFO[98][29] , \FIFO[98][28] ,
         \FIFO[98][27] , \FIFO[98][26] , \FIFO[98][25] , \FIFO[98][24] ,
         \FIFO[98][23] , \FIFO[98][22] , \FIFO[98][21] , \FIFO[98][20] ,
         \FIFO[98][19] , \FIFO[98][18] , \FIFO[98][17] , \FIFO[98][16] ,
         \FIFO[98][15] , \FIFO[98][14] , \FIFO[98][13] , \FIFO[98][12] ,
         \FIFO[98][11] , \FIFO[98][10] , \FIFO[98][9] , \FIFO[98][8] ,
         \FIFO[98][7] , \FIFO[98][6] , \FIFO[98][5] , \FIFO[98][4] ,
         \FIFO[98][3] , \FIFO[98][2] , \FIFO[98][1] , \FIFO[98][0] ,
         \FIFO[99][31] , \FIFO[99][30] , \FIFO[99][29] , \FIFO[99][28] ,
         \FIFO[99][27] , \FIFO[99][26] , \FIFO[99][25] , \FIFO[99][24] ,
         \FIFO[99][23] , \FIFO[99][22] , \FIFO[99][21] , \FIFO[99][20] ,
         \FIFO[99][19] , \FIFO[99][18] , \FIFO[99][17] , \FIFO[99][16] ,
         \FIFO[99][15] , \FIFO[99][14] , \FIFO[99][13] , \FIFO[99][12] ,
         \FIFO[99][11] , \FIFO[99][10] , \FIFO[99][9] , \FIFO[99][8] ,
         \FIFO[99][7] , \FIFO[99][6] , \FIFO[99][5] , \FIFO[99][4] ,
         \FIFO[99][3] , \FIFO[99][2] , \FIFO[99][1] , \FIFO[99][0] ,
         \FIFO[100][31] , \FIFO[100][30] , \FIFO[100][29] , \FIFO[100][28] ,
         \FIFO[100][27] , \FIFO[100][26] , \FIFO[100][25] , \FIFO[100][24] ,
         \FIFO[100][23] , \FIFO[100][22] , \FIFO[100][21] , \FIFO[100][20] ,
         \FIFO[100][19] , \FIFO[100][18] , \FIFO[100][17] , \FIFO[100][16] ,
         \FIFO[100][15] , \FIFO[100][14] , \FIFO[100][13] , \FIFO[100][12] ,
         \FIFO[100][11] , \FIFO[100][10] , \FIFO[100][9] , \FIFO[100][8] ,
         \FIFO[100][7] , \FIFO[100][6] , \FIFO[100][5] , \FIFO[100][4] ,
         \FIFO[100][3] , \FIFO[100][2] , \FIFO[100][1] , \FIFO[100][0] ,
         \FIFO[101][31] , \FIFO[101][30] , \FIFO[101][29] , \FIFO[101][28] ,
         \FIFO[101][27] , \FIFO[101][26] , \FIFO[101][25] , \FIFO[101][24] ,
         \FIFO[101][23] , \FIFO[101][22] , \FIFO[101][21] , \FIFO[101][20] ,
         \FIFO[101][19] , \FIFO[101][18] , \FIFO[101][17] , \FIFO[101][16] ,
         \FIFO[101][15] , \FIFO[101][14] , \FIFO[101][13] , \FIFO[101][12] ,
         \FIFO[101][11] , \FIFO[101][10] , \FIFO[101][9] , \FIFO[101][8] ,
         \FIFO[101][7] , \FIFO[101][6] , \FIFO[101][5] , \FIFO[101][4] ,
         \FIFO[101][3] , \FIFO[101][2] , \FIFO[101][1] , \FIFO[101][0] ,
         \FIFO[102][31] , \FIFO[102][30] , \FIFO[102][29] , \FIFO[102][28] ,
         \FIFO[102][27] , \FIFO[102][26] , \FIFO[102][25] , \FIFO[102][24] ,
         \FIFO[102][23] , \FIFO[102][22] , \FIFO[102][21] , \FIFO[102][20] ,
         \FIFO[102][19] , \FIFO[102][18] , \FIFO[102][17] , \FIFO[102][16] ,
         \FIFO[102][15] , \FIFO[102][14] , \FIFO[102][13] , \FIFO[102][12] ,
         \FIFO[102][11] , \FIFO[102][10] , \FIFO[102][9] , \FIFO[102][8] ,
         \FIFO[102][7] , \FIFO[102][6] , \FIFO[102][5] , \FIFO[102][4] ,
         \FIFO[102][3] , \FIFO[102][2] , \FIFO[102][1] , \FIFO[102][0] ,
         \FIFO[103][31] , \FIFO[103][30] , \FIFO[103][29] , \FIFO[103][28] ,
         \FIFO[103][27] , \FIFO[103][26] , \FIFO[103][25] , \FIFO[103][24] ,
         \FIFO[103][23] , \FIFO[103][22] , \FIFO[103][21] , \FIFO[103][20] ,
         \FIFO[103][19] , \FIFO[103][18] , \FIFO[103][17] , \FIFO[103][16] ,
         \FIFO[103][15] , \FIFO[103][14] , \FIFO[103][13] , \FIFO[103][12] ,
         \FIFO[103][11] , \FIFO[103][10] , \FIFO[103][9] , \FIFO[103][8] ,
         \FIFO[103][7] , \FIFO[103][6] , \FIFO[103][5] , \FIFO[103][4] ,
         \FIFO[103][3] , \FIFO[103][2] , \FIFO[103][1] , \FIFO[103][0] ,
         \FIFO[104][31] , \FIFO[104][30] , \FIFO[104][29] , \FIFO[104][28] ,
         \FIFO[104][27] , \FIFO[104][26] , \FIFO[104][25] , \FIFO[104][24] ,
         \FIFO[104][23] , \FIFO[104][22] , \FIFO[104][21] , \FIFO[104][20] ,
         \FIFO[104][19] , \FIFO[104][18] , \FIFO[104][17] , \FIFO[104][16] ,
         \FIFO[104][15] , \FIFO[104][14] , \FIFO[104][13] , \FIFO[104][12] ,
         \FIFO[104][11] , \FIFO[104][10] , \FIFO[104][9] , \FIFO[104][8] ,
         \FIFO[104][7] , \FIFO[104][6] , \FIFO[104][5] , \FIFO[104][4] ,
         \FIFO[104][3] , \FIFO[104][2] , \FIFO[104][1] , \FIFO[104][0] ,
         \FIFO[105][31] , \FIFO[105][30] , \FIFO[105][29] , \FIFO[105][28] ,
         \FIFO[105][27] , \FIFO[105][26] , \FIFO[105][25] , \FIFO[105][24] ,
         \FIFO[105][23] , \FIFO[105][22] , \FIFO[105][21] , \FIFO[105][20] ,
         \FIFO[105][19] , \FIFO[105][18] , \FIFO[105][17] , \FIFO[105][16] ,
         \FIFO[105][15] , \FIFO[105][14] , \FIFO[105][13] , \FIFO[105][12] ,
         \FIFO[105][11] , \FIFO[105][10] , \FIFO[105][9] , \FIFO[105][8] ,
         \FIFO[105][7] , \FIFO[105][6] , \FIFO[105][5] , \FIFO[105][4] ,
         \FIFO[105][3] , \FIFO[105][2] , \FIFO[105][1] , \FIFO[105][0] ,
         \FIFO[106][31] , \FIFO[106][30] , \FIFO[106][29] , \FIFO[106][28] ,
         \FIFO[106][27] , \FIFO[106][26] , \FIFO[106][25] , \FIFO[106][24] ,
         \FIFO[106][23] , \FIFO[106][22] , \FIFO[106][21] , \FIFO[106][20] ,
         \FIFO[106][19] , \FIFO[106][18] , \FIFO[106][17] , \FIFO[106][16] ,
         \FIFO[106][15] , \FIFO[106][14] , \FIFO[106][13] , \FIFO[106][12] ,
         \FIFO[106][11] , \FIFO[106][10] , \FIFO[106][9] , \FIFO[106][8] ,
         \FIFO[106][7] , \FIFO[106][6] , \FIFO[106][5] , \FIFO[106][4] ,
         \FIFO[106][3] , \FIFO[106][2] , \FIFO[106][1] , \FIFO[106][0] ,
         \FIFO[107][31] , \FIFO[107][30] , \FIFO[107][29] , \FIFO[107][28] ,
         \FIFO[107][27] , \FIFO[107][26] , \FIFO[107][25] , \FIFO[107][24] ,
         \FIFO[107][23] , \FIFO[107][22] , \FIFO[107][21] , \FIFO[107][20] ,
         \FIFO[107][19] , \FIFO[107][18] , \FIFO[107][17] , \FIFO[107][16] ,
         \FIFO[107][15] , \FIFO[107][14] , \FIFO[107][13] , \FIFO[107][12] ,
         \FIFO[107][11] , \FIFO[107][10] , \FIFO[107][9] , \FIFO[107][8] ,
         \FIFO[107][7] , \FIFO[107][6] , \FIFO[107][5] , \FIFO[107][4] ,
         \FIFO[107][3] , \FIFO[107][2] , \FIFO[107][1] , \FIFO[107][0] ,
         \FIFO[108][31] , \FIFO[108][30] , \FIFO[108][29] , \FIFO[108][28] ,
         \FIFO[108][27] , \FIFO[108][26] , \FIFO[108][25] , \FIFO[108][24] ,
         \FIFO[108][23] , \FIFO[108][22] , \FIFO[108][21] , \FIFO[108][20] ,
         \FIFO[108][19] , \FIFO[108][18] , \FIFO[108][17] , \FIFO[108][16] ,
         \FIFO[108][15] , \FIFO[108][14] , \FIFO[108][13] , \FIFO[108][12] ,
         \FIFO[108][11] , \FIFO[108][10] , \FIFO[108][9] , \FIFO[108][8] ,
         \FIFO[108][7] , \FIFO[108][6] , \FIFO[108][5] , \FIFO[108][4] ,
         \FIFO[108][3] , \FIFO[108][2] , \FIFO[108][1] , \FIFO[108][0] ,
         \FIFO[109][31] , \FIFO[109][30] , \FIFO[109][29] , \FIFO[109][28] ,
         \FIFO[109][27] , \FIFO[109][26] , \FIFO[109][25] , \FIFO[109][24] ,
         \FIFO[109][23] , \FIFO[109][22] , \FIFO[109][21] , \FIFO[109][20] ,
         \FIFO[109][19] , \FIFO[109][18] , \FIFO[109][17] , \FIFO[109][16] ,
         \FIFO[109][15] , \FIFO[109][14] , \FIFO[109][13] , \FIFO[109][12] ,
         \FIFO[109][11] , \FIFO[109][10] , \FIFO[109][9] , \FIFO[109][8] ,
         \FIFO[109][7] , \FIFO[109][6] , \FIFO[109][5] , \FIFO[109][4] ,
         \FIFO[109][3] , \FIFO[109][2] , \FIFO[109][1] , \FIFO[109][0] ,
         \FIFO[110][31] , \FIFO[110][30] , \FIFO[110][29] , \FIFO[110][28] ,
         \FIFO[110][27] , \FIFO[110][26] , \FIFO[110][25] , \FIFO[110][24] ,
         \FIFO[110][23] , \FIFO[110][22] , \FIFO[110][21] , \FIFO[110][20] ,
         \FIFO[110][19] , \FIFO[110][18] , \FIFO[110][17] , \FIFO[110][16] ,
         \FIFO[110][15] , \FIFO[110][14] , \FIFO[110][13] , \FIFO[110][12] ,
         \FIFO[110][11] , \FIFO[110][10] , \FIFO[110][9] , \FIFO[110][8] ,
         \FIFO[110][7] , \FIFO[110][6] , \FIFO[110][5] , \FIFO[110][4] ,
         \FIFO[110][3] , \FIFO[110][2] , \FIFO[110][1] , \FIFO[110][0] ,
         \FIFO[111][31] , \FIFO[111][30] , \FIFO[111][29] , \FIFO[111][28] ,
         \FIFO[111][27] , \FIFO[111][26] , \FIFO[111][25] , \FIFO[111][24] ,
         \FIFO[111][23] , \FIFO[111][22] , \FIFO[111][21] , \FIFO[111][20] ,
         \FIFO[111][19] , \FIFO[111][18] , \FIFO[111][17] , \FIFO[111][16] ,
         \FIFO[111][15] , \FIFO[111][14] , \FIFO[111][13] , \FIFO[111][12] ,
         \FIFO[111][11] , \FIFO[111][10] , \FIFO[111][9] , \FIFO[111][8] ,
         \FIFO[111][7] , \FIFO[111][6] , \FIFO[111][5] , \FIFO[111][4] ,
         \FIFO[111][3] , \FIFO[111][2] , \FIFO[111][1] , \FIFO[111][0] ,
         \FIFO[112][31] , \FIFO[112][30] , \FIFO[112][29] , \FIFO[112][28] ,
         \FIFO[112][27] , \FIFO[112][26] , \FIFO[112][25] , \FIFO[112][24] ,
         \FIFO[112][23] , \FIFO[112][22] , \FIFO[112][21] , \FIFO[112][20] ,
         \FIFO[112][19] , \FIFO[112][18] , \FIFO[112][17] , \FIFO[112][16] ,
         \FIFO[112][15] , \FIFO[112][14] , \FIFO[112][13] , \FIFO[112][12] ,
         \FIFO[112][11] , \FIFO[112][10] , \FIFO[112][9] , \FIFO[112][8] ,
         \FIFO[112][7] , \FIFO[112][6] , \FIFO[112][5] , \FIFO[112][4] ,
         \FIFO[112][3] , \FIFO[112][2] , \FIFO[112][1] , \FIFO[112][0] ,
         \FIFO[113][31] , \FIFO[113][30] , \FIFO[113][29] , \FIFO[113][28] ,
         \FIFO[113][27] , \FIFO[113][26] , \FIFO[113][25] , \FIFO[113][24] ,
         \FIFO[113][23] , \FIFO[113][22] , \FIFO[113][21] , \FIFO[113][20] ,
         \FIFO[113][19] , \FIFO[113][18] , \FIFO[113][17] , \FIFO[113][16] ,
         \FIFO[113][15] , \FIFO[113][14] , \FIFO[113][13] , \FIFO[113][12] ,
         \FIFO[113][11] , \FIFO[113][10] , \FIFO[113][9] , \FIFO[113][8] ,
         \FIFO[113][7] , \FIFO[113][6] , \FIFO[113][5] , \FIFO[113][4] ,
         \FIFO[113][3] , \FIFO[113][2] , \FIFO[113][1] , \FIFO[113][0] ,
         \FIFO[114][31] , \FIFO[114][30] , \FIFO[114][29] , \FIFO[114][28] ,
         \FIFO[114][27] , \FIFO[114][26] , \FIFO[114][25] , \FIFO[114][24] ,
         \FIFO[114][23] , \FIFO[114][22] , \FIFO[114][21] , \FIFO[114][20] ,
         \FIFO[114][19] , \FIFO[114][18] , \FIFO[114][17] , \FIFO[114][16] ,
         \FIFO[114][15] , \FIFO[114][14] , \FIFO[114][13] , \FIFO[114][12] ,
         \FIFO[114][11] , \FIFO[114][10] , \FIFO[114][9] , \FIFO[114][8] ,
         \FIFO[114][7] , \FIFO[114][6] , \FIFO[114][5] , \FIFO[114][4] ,
         \FIFO[114][3] , \FIFO[114][2] , \FIFO[114][1] , \FIFO[114][0] ,
         \FIFO[115][31] , \FIFO[115][30] , \FIFO[115][29] , \FIFO[115][28] ,
         \FIFO[115][27] , \FIFO[115][26] , \FIFO[115][25] , \FIFO[115][24] ,
         \FIFO[115][23] , \FIFO[115][22] , \FIFO[115][21] , \FIFO[115][20] ,
         \FIFO[115][19] , \FIFO[115][18] , \FIFO[115][17] , \FIFO[115][16] ,
         \FIFO[115][15] , \FIFO[115][14] , \FIFO[115][13] , \FIFO[115][12] ,
         \FIFO[115][11] , \FIFO[115][10] , \FIFO[115][9] , \FIFO[115][8] ,
         \FIFO[115][7] , \FIFO[115][6] , \FIFO[115][5] , \FIFO[115][4] ,
         \FIFO[115][3] , \FIFO[115][2] , \FIFO[115][1] , \FIFO[115][0] ,
         \FIFO[116][31] , \FIFO[116][30] , \FIFO[116][29] , \FIFO[116][28] ,
         \FIFO[116][27] , \FIFO[116][26] , \FIFO[116][25] , \FIFO[116][24] ,
         \FIFO[116][23] , \FIFO[116][22] , \FIFO[116][21] , \FIFO[116][20] ,
         \FIFO[116][19] , \FIFO[116][18] , \FIFO[116][17] , \FIFO[116][16] ,
         \FIFO[116][15] , \FIFO[116][14] , \FIFO[116][13] , \FIFO[116][12] ,
         \FIFO[116][11] , \FIFO[116][10] , \FIFO[116][9] , \FIFO[116][8] ,
         \FIFO[116][7] , \FIFO[116][6] , \FIFO[116][5] , \FIFO[116][4] ,
         \FIFO[116][3] , \FIFO[116][2] , \FIFO[116][1] , \FIFO[116][0] ,
         \FIFO[117][31] , \FIFO[117][30] , \FIFO[117][29] , \FIFO[117][28] ,
         \FIFO[117][27] , \FIFO[117][26] , \FIFO[117][25] , \FIFO[117][24] ,
         \FIFO[117][23] , \FIFO[117][22] , \FIFO[117][21] , \FIFO[117][20] ,
         \FIFO[117][19] , \FIFO[117][18] , \FIFO[117][17] , \FIFO[117][16] ,
         \FIFO[117][15] , \FIFO[117][14] , \FIFO[117][13] , \FIFO[117][12] ,
         \FIFO[117][11] , \FIFO[117][10] , \FIFO[117][9] , \FIFO[117][8] ,
         \FIFO[117][7] , \FIFO[117][6] , \FIFO[117][5] , \FIFO[117][4] ,
         \FIFO[117][3] , \FIFO[117][2] , \FIFO[117][1] , \FIFO[117][0] ,
         \FIFO[118][31] , \FIFO[118][30] , \FIFO[118][29] , \FIFO[118][28] ,
         \FIFO[118][27] , \FIFO[118][26] , \FIFO[118][25] , \FIFO[118][24] ,
         \FIFO[118][23] , \FIFO[118][22] , \FIFO[118][21] , \FIFO[118][20] ,
         \FIFO[118][19] , \FIFO[118][18] , \FIFO[118][17] , \FIFO[118][16] ,
         \FIFO[118][15] , \FIFO[118][14] , \FIFO[118][13] , \FIFO[118][12] ,
         \FIFO[118][11] , \FIFO[118][10] , \FIFO[118][9] , \FIFO[118][8] ,
         \FIFO[118][7] , \FIFO[118][6] , \FIFO[118][5] , \FIFO[118][4] ,
         \FIFO[118][3] , \FIFO[118][2] , \FIFO[118][1] , \FIFO[118][0] ,
         \FIFO[119][31] , \FIFO[119][30] , \FIFO[119][29] , \FIFO[119][28] ,
         \FIFO[119][27] , \FIFO[119][26] , \FIFO[119][25] , \FIFO[119][24] ,
         \FIFO[119][23] , \FIFO[119][22] , \FIFO[119][21] , \FIFO[119][20] ,
         \FIFO[119][19] , \FIFO[119][18] , \FIFO[119][17] , \FIFO[119][16] ,
         \FIFO[119][15] , \FIFO[119][14] , \FIFO[119][13] , \FIFO[119][12] ,
         \FIFO[119][11] , \FIFO[119][10] , \FIFO[119][9] , \FIFO[119][8] ,
         \FIFO[119][7] , \FIFO[119][6] , \FIFO[119][5] , \FIFO[119][4] ,
         \FIFO[119][3] , \FIFO[119][2] , \FIFO[119][1] , \FIFO[119][0] ,
         \FIFO[120][31] , \FIFO[120][30] , \FIFO[120][29] , \FIFO[120][28] ,
         \FIFO[120][27] , \FIFO[120][26] , \FIFO[120][25] , \FIFO[120][24] ,
         \FIFO[120][23] , \FIFO[120][22] , \FIFO[120][21] , \FIFO[120][20] ,
         \FIFO[120][19] , \FIFO[120][18] , \FIFO[120][17] , \FIFO[120][16] ,
         \FIFO[120][15] , \FIFO[120][14] , \FIFO[120][13] , \FIFO[120][12] ,
         \FIFO[120][11] , \FIFO[120][10] , \FIFO[120][9] , \FIFO[120][8] ,
         \FIFO[120][7] , \FIFO[120][6] , \FIFO[120][5] , \FIFO[120][4] ,
         \FIFO[120][3] , \FIFO[120][2] , \FIFO[120][1] , \FIFO[120][0] ,
         \FIFO[121][31] , \FIFO[121][30] , \FIFO[121][29] , \FIFO[121][28] ,
         \FIFO[121][27] , \FIFO[121][26] , \FIFO[121][25] , \FIFO[121][24] ,
         \FIFO[121][23] , \FIFO[121][22] , \FIFO[121][21] , \FIFO[121][20] ,
         \FIFO[121][19] , \FIFO[121][18] , \FIFO[121][17] , \FIFO[121][16] ,
         \FIFO[121][15] , \FIFO[121][14] , \FIFO[121][13] , \FIFO[121][12] ,
         \FIFO[121][11] , \FIFO[121][10] , \FIFO[121][9] , \FIFO[121][8] ,
         \FIFO[121][7] , \FIFO[121][6] , \FIFO[121][5] , \FIFO[121][4] ,
         \FIFO[121][3] , \FIFO[121][2] , \FIFO[121][1] , \FIFO[121][0] ,
         \FIFO[122][31] , \FIFO[122][30] , \FIFO[122][29] , \FIFO[122][28] ,
         \FIFO[122][27] , \FIFO[122][26] , \FIFO[122][25] , \FIFO[122][24] ,
         \FIFO[122][23] , \FIFO[122][22] , \FIFO[122][21] , \FIFO[122][20] ,
         \FIFO[122][19] , \FIFO[122][18] , \FIFO[122][17] , \FIFO[122][16] ,
         \FIFO[122][15] , \FIFO[122][14] , \FIFO[122][13] , \FIFO[122][12] ,
         \FIFO[122][11] , \FIFO[122][10] , \FIFO[122][9] , \FIFO[122][8] ,
         \FIFO[122][7] , \FIFO[122][6] , \FIFO[122][5] , \FIFO[122][4] ,
         \FIFO[122][3] , \FIFO[122][2] , \FIFO[122][1] , \FIFO[122][0] ,
         \FIFO[123][31] , \FIFO[123][30] , \FIFO[123][29] , \FIFO[123][28] ,
         \FIFO[123][27] , \FIFO[123][26] , \FIFO[123][25] , \FIFO[123][24] ,
         \FIFO[123][23] , \FIFO[123][22] , \FIFO[123][21] , \FIFO[123][20] ,
         \FIFO[123][19] , \FIFO[123][18] , \FIFO[123][17] , \FIFO[123][16] ,
         \FIFO[123][15] , \FIFO[123][14] , \FIFO[123][13] , \FIFO[123][12] ,
         \FIFO[123][11] , \FIFO[123][10] , \FIFO[123][9] , \FIFO[123][8] ,
         \FIFO[123][7] , \FIFO[123][6] , \FIFO[123][5] , \FIFO[123][4] ,
         \FIFO[123][3] , \FIFO[123][2] , \FIFO[123][1] , \FIFO[123][0] ,
         \FIFO[124][31] , \FIFO[124][30] , \FIFO[124][29] , \FIFO[124][28] ,
         \FIFO[124][27] , \FIFO[124][26] , \FIFO[124][25] , \FIFO[124][24] ,
         \FIFO[124][23] , \FIFO[124][22] , \FIFO[124][21] , \FIFO[124][20] ,
         \FIFO[124][19] , \FIFO[124][18] , \FIFO[124][17] , \FIFO[124][16] ,
         \FIFO[124][15] , \FIFO[124][14] , \FIFO[124][13] , \FIFO[124][12] ,
         \FIFO[124][11] , \FIFO[124][10] , \FIFO[124][9] , \FIFO[124][8] ,
         \FIFO[124][7] , \FIFO[124][6] , \FIFO[124][5] , \FIFO[124][4] ,
         \FIFO[124][3] , \FIFO[124][2] , \FIFO[124][1] , \FIFO[124][0] ,
         \FIFO[125][31] , \FIFO[125][30] , \FIFO[125][29] , \FIFO[125][28] ,
         \FIFO[125][27] , \FIFO[125][26] , \FIFO[125][25] , \FIFO[125][24] ,
         \FIFO[125][23] , \FIFO[125][22] , \FIFO[125][21] , \FIFO[125][20] ,
         \FIFO[125][19] , \FIFO[125][18] , \FIFO[125][17] , \FIFO[125][16] ,
         \FIFO[125][15] , \FIFO[125][14] , \FIFO[125][13] , \FIFO[125][12] ,
         \FIFO[125][11] , \FIFO[125][10] , \FIFO[125][9] , \FIFO[125][8] ,
         \FIFO[125][7] , \FIFO[125][6] , \FIFO[125][5] , \FIFO[125][4] ,
         \FIFO[125][3] , \FIFO[125][2] , \FIFO[125][1] , \FIFO[125][0] ,
         \FIFO[126][31] , \FIFO[126][30] , \FIFO[126][29] , \FIFO[126][28] ,
         \FIFO[126][27] , \FIFO[126][26] , \FIFO[126][25] , \FIFO[126][24] ,
         \FIFO[126][23] , \FIFO[126][22] , \FIFO[126][21] , \FIFO[126][20] ,
         \FIFO[126][19] , \FIFO[126][18] , \FIFO[126][17] , \FIFO[126][16] ,
         \FIFO[126][15] , \FIFO[126][14] , \FIFO[126][13] , \FIFO[126][12] ,
         \FIFO[126][11] , \FIFO[126][10] , \FIFO[126][9] , \FIFO[126][8] ,
         \FIFO[126][7] , \FIFO[126][6] , \FIFO[126][5] , \FIFO[126][4] ,
         \FIFO[126][3] , \FIFO[126][2] , \FIFO[126][1] , \FIFO[126][0] ,
         \FIFO[127][31] , \FIFO[127][30] , \FIFO[127][29] , \FIFO[127][28] ,
         \FIFO[127][27] , \FIFO[127][26] , \FIFO[127][25] , \FIFO[127][24] ,
         \FIFO[127][23] , \FIFO[127][22] , \FIFO[127][21] , \FIFO[127][20] ,
         \FIFO[127][19] , \FIFO[127][18] , \FIFO[127][17] , \FIFO[127][16] ,
         \FIFO[127][15] , \FIFO[127][14] , \FIFO[127][13] , \FIFO[127][12] ,
         \FIFO[127][11] , \FIFO[127][10] , \FIFO[127][9] , \FIFO[127][8] ,
         \FIFO[127][7] , \FIFO[127][6] , \FIFO[127][5] , \FIFO[127][4] ,
         \FIFO[127][3] , \FIFO[127][2] , \FIFO[127][1] , \FIFO[127][0] , N219,
         N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230,
         N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241,
         N242, N243, N244, N245, N246, N247, N248, N249, N250, N253, N254,
         N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, N265,
         N266, N267, N268, N269, N270, N271, N272, N273, N274, N275, N276,
         N277, N278, N279, N280, N281, N282, N283, n204, n206, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n400, n401, n464, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n205, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n398, n399, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n465, n466, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368;
  assign N15 = rdaddr[0];
  assign N16 = rdaddr[1];
  assign N17 = rdaddr[2];
  assign N18 = rdaddr[3];
  assign N19 = rdaddr[4];
  assign N20 = rdaddr[5];
  assign N21 = rdaddr[6];
  assign sync_flush = sync_flush_BAR;
  assign wren = wren_BAR;

  DFFARX1 \FIFO_reg[0][31]  ( .D(n4562), .CLK(clk_in), .RSTB(n7106), .Q(
        \FIFO[0][31] ), .QN(n19) );
  DFFARX1 \FIFO_reg[0][30]  ( .D(n4561), .CLK(clk_in), .RSTB(n7106), .Q(
        \FIFO[0][30] ), .QN(n15) );
  DFFARX1 \FIFO_reg[0][29]  ( .D(n4560), .CLK(clk_in), .RSTB(n7106), .Q(
        \FIFO[0][29] ), .QN(n13) );
  DFFARX1 \FIFO_reg[0][28]  ( .D(n4559), .CLK(clk_in), .RSTB(n7106), .Q(
        \FIFO[0][28] ) );
  DFFARX1 \FIFO_reg[0][27]  ( .D(n4558), .CLK(clk_in), .RSTB(n7106), .Q(
        \FIFO[0][27] ), .QN(n10) );
  DFFARX1 \FIFO_reg[0][26]  ( .D(n4557), .CLK(clk_in), .RSTB(n7106), .Q(
        \FIFO[0][26] ) );
  DFFARX1 \FIFO_reg[0][25]  ( .D(n4556), .CLK(clk_in), .RSTB(n7107), .Q(
        \FIFO[0][25] ) );
  DFFARX1 \FIFO_reg[0][24]  ( .D(n4555), .CLK(clk_in), .RSTB(n7107), .Q(
        \FIFO[0][24] ) );
  DFFARX1 \FIFO_reg[0][23]  ( .D(n4554), .CLK(clk_in), .RSTB(n7107), .Q(
        \FIFO[0][23] ), .QN(n16) );
  DFFARX1 \FIFO_reg[0][22]  ( .D(n4553), .CLK(clk_in), .RSTB(n7107), .Q(
        \FIFO[0][22] ), .QN(n18) );
  DFFARX1 \FIFO_reg[0][21]  ( .D(n4552), .CLK(clk_in), .RSTB(n7107), .Q(
        \FIFO[0][21] ), .QN(n12) );
  DFFARX1 \FIFO_reg[0][20]  ( .D(n4551), .CLK(clk_in), .RSTB(n7107), .Q(
        \FIFO[0][20] ), .QN(n9) );
  DFFARX1 \FIFO_reg[0][19]  ( .D(n4550), .CLK(clk_in), .RSTB(n7107), .Q(
        \FIFO[0][19] ) );
  DFFARX1 \FIFO_reg[0][18]  ( .D(n4549), .CLK(clk_in), .RSTB(n7107), .Q(
        \FIFO[0][18] ) );
  DFFARX1 \FIFO_reg[0][17]  ( .D(n4548), .CLK(clk_in), .RSTB(n7107), .Q(
        \FIFO[0][17] ) );
  DFFARX1 \FIFO_reg[0][16]  ( .D(n4547), .CLK(clk_in), .RSTB(n7107), .Q(
        \FIFO[0][16] ) );
  DFFARX1 \FIFO_reg[0][15]  ( .D(n4546), .CLK(clk_in), .RSTB(n7107), .Q(
        \FIFO[0][15] ) );
  DFFARX1 \FIFO_reg[0][14]  ( .D(n4545), .CLK(clk_in), .RSTB(n7107), .Q(
        \FIFO[0][14] ) );
  DFFARX1 \FIFO_reg[0][13]  ( .D(n4544), .CLK(clk_in), .RSTB(n7107), .Q(
        \FIFO[0][13] ) );
  DFFARX1 \FIFO_reg[0][12]  ( .D(n4543), .CLK(clk_in), .RSTB(n7107), .Q(
        \FIFO[0][12] ) );
  DFFARX1 \FIFO_reg[0][11]  ( .D(n4542), .CLK(clk_in), .RSTB(n7107), .Q(
        \FIFO[0][11] ), .QN(n17) );
  DFFARX1 \FIFO_reg[0][10]  ( .D(n4541), .CLK(clk_in), .RSTB(n7107), .Q(
        \FIFO[0][10] ), .QN(n14) );
  DFFARX1 \FIFO_reg[0][9]  ( .D(n4540), .CLK(clk_in), .RSTB(n7107), .Q(
        \FIFO[0][9] ), .QN(n11) );
  DFFARX1 \FIFO_reg[0][8]  ( .D(n4539), .CLK(clk_in), .RSTB(n7107), .Q(
        \FIFO[0][8] ) );
  DFFARX1 \FIFO_reg[0][7]  ( .D(n4538), .CLK(clk_in), .RSTB(n7108), .Q(
        \FIFO[0][7] ) );
  DFFARX1 \FIFO_reg[0][6]  ( .D(n4537), .CLK(clk_in), .RSTB(n7108), .Q(
        \FIFO[0][6] ) );
  DFFARX1 \FIFO_reg[0][5]  ( .D(n4536), .CLK(clk_in), .RSTB(n7108), .Q(
        \FIFO[0][5] ) );
  DFFARX1 \FIFO_reg[0][4]  ( .D(n4535), .CLK(clk_in), .RSTB(n7108), .Q(
        \FIFO[0][4] ) );
  DFFARX1 \FIFO_reg[0][3]  ( .D(n4534), .CLK(clk_in), .RSTB(n7108), .Q(
        \FIFO[0][3] ) );
  DFFARX1 \FIFO_reg[0][2]  ( .D(n4533), .CLK(clk_in), .RSTB(n7108), .Q(
        \FIFO[0][2] ) );
  DFFARX1 \FIFO_reg[0][1]  ( .D(n4532), .CLK(clk_in), .RSTB(n7108), .Q(
        \FIFO[0][1] ) );
  DFFARX1 \FIFO_reg[0][0]  ( .D(n4531), .CLK(clk_in), .RSTB(n7108), .Q(
        \FIFO[0][0] ) );
  DFFARX1 \FIFO_reg[1][31]  ( .D(n4530), .CLK(clk_in), .RSTB(n7108), .Q(
        \FIFO[1][31] ) );
  DFFARX1 \FIFO_reg[1][30]  ( .D(n4529), .CLK(clk_in), .RSTB(n7108), .Q(
        \FIFO[1][30] ) );
  DFFARX1 \FIFO_reg[1][29]  ( .D(n4528), .CLK(clk_in), .RSTB(n7108), .Q(
        \FIFO[1][29] ) );
  DFFARX1 \FIFO_reg[1][28]  ( .D(n4527), .CLK(clk_in), .RSTB(n7108), .Q(
        \FIFO[1][28] ) );
  DFFARX1 \FIFO_reg[1][27]  ( .D(n4526), .CLK(clk_in), .RSTB(n7108), .Q(
        \FIFO[1][27] ) );
  DFFARX1 \FIFO_reg[1][26]  ( .D(n4525), .CLK(clk_in), .RSTB(n7108), .Q(
        \FIFO[1][26] ) );
  DFFARX1 \FIFO_reg[1][25]  ( .D(n4524), .CLK(clk_in), .RSTB(n7108), .Q(
        \FIFO[1][25] ) );
  DFFARX1 \FIFO_reg[1][24]  ( .D(n4523), .CLK(clk_in), .RSTB(n7108), .Q(
        \FIFO[1][24] ) );
  DFFARX1 \FIFO_reg[1][23]  ( .D(n4522), .CLK(clk_in), .RSTB(n7108), .Q(
        \FIFO[1][23] ) );
  DFFARX1 \FIFO_reg[1][22]  ( .D(n4521), .CLK(clk_in), .RSTB(n7108), .Q(
        \FIFO[1][22] ) );
  DFFARX1 \FIFO_reg[1][21]  ( .D(n4520), .CLK(clk_in), .RSTB(n7109), .Q(
        \FIFO[1][21] ) );
  DFFARX1 \FIFO_reg[1][20]  ( .D(n4519), .CLK(clk_in), .RSTB(n7109), .Q(
        \FIFO[1][20] ) );
  DFFARX1 \FIFO_reg[1][19]  ( .D(n4518), .CLK(clk_in), .RSTB(n7109), .Q(
        \FIFO[1][19] ) );
  DFFARX1 \FIFO_reg[1][18]  ( .D(n4517), .CLK(clk_in), .RSTB(n7109), .Q(
        \FIFO[1][18] ) );
  DFFARX1 \FIFO_reg[1][17]  ( .D(n4516), .CLK(clk_in), .RSTB(n7109), .Q(
        \FIFO[1][17] ) );
  DFFARX1 \FIFO_reg[1][16]  ( .D(n4515), .CLK(clk_in), .RSTB(n7109), .Q(
        \FIFO[1][16] ) );
  DFFARX1 \FIFO_reg[1][15]  ( .D(n4514), .CLK(clk_in), .RSTB(n7109), .Q(
        \FIFO[1][15] ) );
  DFFARX1 \FIFO_reg[1][14]  ( .D(n4513), .CLK(clk_in), .RSTB(n7109), .Q(
        \FIFO[1][14] ) );
  DFFARX1 \FIFO_reg[1][13]  ( .D(n4512), .CLK(clk_in), .RSTB(n7109), .Q(
        \FIFO[1][13] ) );
  DFFARX1 \FIFO_reg[1][12]  ( .D(n4511), .CLK(clk_in), .RSTB(n7109), .Q(
        \FIFO[1][12] ) );
  DFFARX1 \FIFO_reg[1][11]  ( .D(n4510), .CLK(clk_in), .RSTB(n7109), .Q(
        \FIFO[1][11] ) );
  DFFARX1 \FIFO_reg[1][10]  ( .D(n4509), .CLK(clk_in), .RSTB(n7109), .Q(
        \FIFO[1][10] ) );
  DFFARX1 \FIFO_reg[1][9]  ( .D(n4508), .CLK(clk_in), .RSTB(n7109), .Q(
        \FIFO[1][9] ) );
  DFFARX1 \FIFO_reg[1][8]  ( .D(n4507), .CLK(clk_in), .RSTB(n7109), .Q(
        \FIFO[1][8] ) );
  DFFARX1 \FIFO_reg[1][7]  ( .D(n4506), .CLK(clk_in), .RSTB(n7109), .Q(
        \FIFO[1][7] ) );
  DFFARX1 \FIFO_reg[1][6]  ( .D(n4505), .CLK(clk_in), .RSTB(n7109), .Q(
        \FIFO[1][6] ) );
  DFFARX1 \FIFO_reg[1][5]  ( .D(n4504), .CLK(clk_in), .RSTB(n7109), .Q(
        \FIFO[1][5] ) );
  DFFARX1 \FIFO_reg[1][4]  ( .D(n4503), .CLK(clk_in), .RSTB(n7109), .Q(
        \FIFO[1][4] ) );
  DFFARX1 \FIFO_reg[1][3]  ( .D(n4502), .CLK(clk_in), .RSTB(n7110), .Q(
        \FIFO[1][3] ) );
  DFFARX1 \FIFO_reg[1][2]  ( .D(n4501), .CLK(clk_in), .RSTB(n7110), .Q(
        \FIFO[1][2] ) );
  DFFARX1 \FIFO_reg[1][1]  ( .D(n4500), .CLK(clk_in), .RSTB(n7110), .Q(
        \FIFO[1][1] ) );
  DFFARX1 \FIFO_reg[1][0]  ( .D(n4499), .CLK(clk_in), .RSTB(n7110), .Q(
        \FIFO[1][0] ) );
  DFFARX1 \FIFO_reg[2][31]  ( .D(n4498), .CLK(clk_in), .RSTB(n7110), .Q(
        \FIFO[2][31] ) );
  DFFARX1 \FIFO_reg[2][30]  ( .D(n4497), .CLK(clk_in), .RSTB(n7110), .Q(
        \FIFO[2][30] ) );
  DFFARX1 \FIFO_reg[2][29]  ( .D(n4496), .CLK(clk_in), .RSTB(n7110), .Q(
        \FIFO[2][29] ) );
  DFFARX1 \FIFO_reg[2][28]  ( .D(n4495), .CLK(clk_in), .RSTB(n7110), .Q(
        \FIFO[2][28] ) );
  DFFARX1 \FIFO_reg[2][27]  ( .D(n4494), .CLK(clk_in), .RSTB(n7110), .Q(
        \FIFO[2][27] ) );
  DFFARX1 \FIFO_reg[2][26]  ( .D(n4493), .CLK(clk_in), .RSTB(n7110), .Q(
        \FIFO[2][26] ) );
  DFFARX1 \FIFO_reg[2][25]  ( .D(n4492), .CLK(clk_in), .RSTB(n7110), .Q(
        \FIFO[2][25] ) );
  DFFARX1 \FIFO_reg[2][24]  ( .D(n4491), .CLK(clk_in), .RSTB(n7110), .Q(
        \FIFO[2][24] ) );
  DFFARX1 \FIFO_reg[2][23]  ( .D(n4490), .CLK(clk_in), .RSTB(n7110), .Q(
        \FIFO[2][23] ) );
  DFFARX1 \FIFO_reg[2][22]  ( .D(n4489), .CLK(clk_in), .RSTB(n7110), .Q(
        \FIFO[2][22] ) );
  DFFARX1 \FIFO_reg[2][21]  ( .D(n4488), .CLK(clk_in), .RSTB(n7110), .Q(
        \FIFO[2][21] ) );
  DFFARX1 \FIFO_reg[2][20]  ( .D(n4487), .CLK(clk_in), .RSTB(n7110), .Q(
        \FIFO[2][20] ) );
  DFFARX1 \FIFO_reg[2][19]  ( .D(n4486), .CLK(clk_in), .RSTB(n7110), .Q(
        \FIFO[2][19] ) );
  DFFARX1 \FIFO_reg[2][18]  ( .D(n4485), .CLK(clk_in), .RSTB(n7110), .Q(
        \FIFO[2][18] ) );
  DFFARX1 \FIFO_reg[2][17]  ( .D(n4484), .CLK(clk_in), .RSTB(n7111), .Q(
        \FIFO[2][17] ) );
  DFFARX1 \FIFO_reg[2][16]  ( .D(n4483), .CLK(clk_in), .RSTB(n7111), .Q(
        \FIFO[2][16] ) );
  DFFARX1 \FIFO_reg[2][15]  ( .D(n4482), .CLK(clk_in), .RSTB(n7111), .Q(
        \FIFO[2][15] ) );
  DFFARX1 \FIFO_reg[2][14]  ( .D(n4481), .CLK(clk_in), .RSTB(n7111), .Q(
        \FIFO[2][14] ) );
  DFFARX1 \FIFO_reg[2][13]  ( .D(n4480), .CLK(clk_in), .RSTB(n7111), .Q(
        \FIFO[2][13] ) );
  DFFARX1 \FIFO_reg[2][12]  ( .D(n4479), .CLK(clk_in), .RSTB(n7111), .Q(
        \FIFO[2][12] ) );
  DFFARX1 \FIFO_reg[2][11]  ( .D(n4478), .CLK(clk_in), .RSTB(n7111), .Q(
        \FIFO[2][11] ) );
  DFFARX1 \FIFO_reg[2][10]  ( .D(n4477), .CLK(clk_in), .RSTB(n7111), .Q(
        \FIFO[2][10] ) );
  DFFARX1 \FIFO_reg[2][9]  ( .D(n4476), .CLK(clk_in), .RSTB(n7111), .Q(
        \FIFO[2][9] ) );
  DFFARX1 \FIFO_reg[2][8]  ( .D(n4475), .CLK(clk_in), .RSTB(n7111), .Q(
        \FIFO[2][8] ) );
  DFFARX1 \FIFO_reg[2][7]  ( .D(n4474), .CLK(clk_in), .RSTB(n7111), .Q(
        \FIFO[2][7] ) );
  DFFARX1 \FIFO_reg[2][6]  ( .D(n4473), .CLK(clk_in), .RSTB(n7111), .Q(
        \FIFO[2][6] ) );
  DFFARX1 \FIFO_reg[2][5]  ( .D(n4472), .CLK(clk_in), .RSTB(n7111), .Q(
        \FIFO[2][5] ) );
  DFFARX1 \FIFO_reg[2][4]  ( .D(n4471), .CLK(clk_in), .RSTB(n7111), .Q(
        \FIFO[2][4] ) );
  DFFARX1 \FIFO_reg[2][3]  ( .D(n4470), .CLK(clk_in), .RSTB(n7111), .Q(
        \FIFO[2][3] ) );
  DFFARX1 \FIFO_reg[2][2]  ( .D(n4469), .CLK(clk_in), .RSTB(n7111), .Q(
        \FIFO[2][2] ) );
  DFFARX1 \FIFO_reg[2][1]  ( .D(n4468), .CLK(clk_in), .RSTB(n7111), .Q(
        \FIFO[2][1] ) );
  DFFARX1 \FIFO_reg[2][0]  ( .D(n4467), .CLK(clk_in), .RSTB(n7111), .Q(
        \FIFO[2][0] ) );
  DFFARX1 \FIFO_reg[3][31]  ( .D(n4466), .CLK(clk_in), .RSTB(n7112), .Q(
        \FIFO[3][31] ) );
  DFFARX1 \FIFO_reg[3][30]  ( .D(n4465), .CLK(clk_in), .RSTB(n7112), .Q(
        \FIFO[3][30] ) );
  DFFARX1 \FIFO_reg[3][29]  ( .D(n4464), .CLK(clk_in), .RSTB(n7112), .Q(
        \FIFO[3][29] ) );
  DFFARX1 \FIFO_reg[3][28]  ( .D(n4463), .CLK(clk_in), .RSTB(n7112), .Q(
        \FIFO[3][28] ) );
  DFFARX1 \FIFO_reg[3][27]  ( .D(n4462), .CLK(clk_in), .RSTB(n7112), .Q(
        \FIFO[3][27] ) );
  DFFARX1 \FIFO_reg[3][26]  ( .D(n4461), .CLK(clk_in), .RSTB(n7112), .Q(
        \FIFO[3][26] ) );
  DFFARX1 \FIFO_reg[3][25]  ( .D(n4460), .CLK(clk_in), .RSTB(n7112), .Q(
        \FIFO[3][25] ) );
  DFFARX1 \FIFO_reg[3][24]  ( .D(n4459), .CLK(clk_in), .RSTB(n7112), .Q(
        \FIFO[3][24] ) );
  DFFARX1 \FIFO_reg[3][23]  ( .D(n4458), .CLK(clk_in), .RSTB(n7112), .Q(
        \FIFO[3][23] ) );
  DFFARX1 \FIFO_reg[3][22]  ( .D(n4457), .CLK(clk_in), .RSTB(n7112), .Q(
        \FIFO[3][22] ) );
  DFFARX1 \FIFO_reg[3][21]  ( .D(n4456), .CLK(clk_in), .RSTB(n7112), .Q(
        \FIFO[3][21] ) );
  DFFARX1 \FIFO_reg[3][20]  ( .D(n4455), .CLK(clk_in), .RSTB(n7112), .Q(
        \FIFO[3][20] ) );
  DFFARX1 \FIFO_reg[3][19]  ( .D(n4454), .CLK(clk_in), .RSTB(n7112), .Q(
        \FIFO[3][19] ) );
  DFFARX1 \FIFO_reg[3][18]  ( .D(n4453), .CLK(clk_in), .RSTB(n7112), .Q(
        \FIFO[3][18] ) );
  DFFARX1 \FIFO_reg[3][17]  ( .D(n4452), .CLK(clk_in), .RSTB(n7112), .Q(
        \FIFO[3][17] ) );
  DFFARX1 \FIFO_reg[3][16]  ( .D(n4451), .CLK(clk_in), .RSTB(n7112), .Q(
        \FIFO[3][16] ) );
  DFFARX1 \FIFO_reg[3][15]  ( .D(n4450), .CLK(clk_in), .RSTB(n7112), .Q(
        \FIFO[3][15] ) );
  DFFARX1 \FIFO_reg[3][14]  ( .D(n4449), .CLK(clk_in), .RSTB(n7112), .Q(
        \FIFO[3][14] ) );
  DFFARX1 \FIFO_reg[3][13]  ( .D(n4448), .CLK(clk_in), .RSTB(n7113), .Q(
        \FIFO[3][13] ) );
  DFFARX1 \FIFO_reg[3][12]  ( .D(n4447), .CLK(clk_in), .RSTB(n7113), .Q(
        \FIFO[3][12] ) );
  DFFARX1 \FIFO_reg[3][11]  ( .D(n4446), .CLK(clk_in), .RSTB(n7113), .Q(
        \FIFO[3][11] ) );
  DFFARX1 \FIFO_reg[3][10]  ( .D(n4445), .CLK(clk_in), .RSTB(n7113), .Q(
        \FIFO[3][10] ) );
  DFFARX1 \FIFO_reg[3][9]  ( .D(n4444), .CLK(clk_in), .RSTB(n7113), .Q(
        \FIFO[3][9] ) );
  DFFARX1 \FIFO_reg[3][8]  ( .D(n4443), .CLK(clk_in), .RSTB(n7113), .Q(
        \FIFO[3][8] ) );
  DFFARX1 \FIFO_reg[3][7]  ( .D(n4442), .CLK(clk_in), .RSTB(n7113), .Q(
        \FIFO[3][7] ) );
  DFFARX1 \FIFO_reg[3][6]  ( .D(n4441), .CLK(clk_in), .RSTB(n7113), .Q(
        \FIFO[3][6] ) );
  DFFARX1 \FIFO_reg[3][5]  ( .D(n4440), .CLK(clk_in), .RSTB(n7113), .Q(
        \FIFO[3][5] ) );
  DFFARX1 \FIFO_reg[3][4]  ( .D(n4439), .CLK(clk_in), .RSTB(n7113), .Q(
        \FIFO[3][4] ) );
  DFFARX1 \FIFO_reg[3][3]  ( .D(n4438), .CLK(clk_in), .RSTB(n7113), .Q(
        \FIFO[3][3] ) );
  DFFARX1 \FIFO_reg[3][2]  ( .D(n4437), .CLK(clk_in), .RSTB(n7113), .Q(
        \FIFO[3][2] ) );
  DFFARX1 \FIFO_reg[3][1]  ( .D(n4436), .CLK(clk_in), .RSTB(n7113), .Q(
        \FIFO[3][1] ) );
  DFFARX1 \FIFO_reg[3][0]  ( .D(n4435), .CLK(clk_in), .RSTB(n7113), .Q(
        \FIFO[3][0] ) );
  DFFARX1 \FIFO_reg[4][31]  ( .D(n4434), .CLK(clk_in), .RSTB(n7113), .Q(
        \FIFO[4][31] ) );
  DFFARX1 \FIFO_reg[4][30]  ( .D(n4433), .CLK(clk_in), .RSTB(n7113), .Q(
        \FIFO[4][30] ) );
  DFFARX1 \FIFO_reg[4][29]  ( .D(n4432), .CLK(clk_in), .RSTB(n7113), .Q(
        \FIFO[4][29] ) );
  DFFARX1 \FIFO_reg[4][28]  ( .D(n4431), .CLK(clk_in), .RSTB(n7113), .Q(
        \FIFO[4][28] ) );
  DFFARX1 \FIFO_reg[4][27]  ( .D(n4430), .CLK(clk_in), .RSTB(n7114), .Q(
        \FIFO[4][27] ) );
  DFFARX1 \FIFO_reg[4][26]  ( .D(n4429), .CLK(clk_in), .RSTB(n7114), .Q(
        \FIFO[4][26] ) );
  DFFARX1 \FIFO_reg[4][25]  ( .D(n4428), .CLK(clk_in), .RSTB(n7114), .Q(
        \FIFO[4][25] ) );
  DFFARX1 \FIFO_reg[4][24]  ( .D(n4427), .CLK(clk_in), .RSTB(n7114), .Q(
        \FIFO[4][24] ) );
  DFFARX1 \FIFO_reg[4][23]  ( .D(n4426), .CLK(clk_in), .RSTB(n7114), .Q(
        \FIFO[4][23] ) );
  DFFARX1 \FIFO_reg[4][22]  ( .D(n4425), .CLK(clk_in), .RSTB(n7114), .Q(
        \FIFO[4][22] ) );
  DFFARX1 \FIFO_reg[4][21]  ( .D(n4424), .CLK(clk_in), .RSTB(n7114), .Q(
        \FIFO[4][21] ) );
  DFFARX1 \FIFO_reg[4][20]  ( .D(n4423), .CLK(clk_in), .RSTB(n7114), .Q(
        \FIFO[4][20] ) );
  DFFARX1 \FIFO_reg[4][19]  ( .D(n4422), .CLK(clk_in), .RSTB(n7114), .Q(
        \FIFO[4][19] ) );
  DFFARX1 \FIFO_reg[4][18]  ( .D(n4421), .CLK(clk_in), .RSTB(n7114), .Q(
        \FIFO[4][18] ) );
  DFFARX1 \FIFO_reg[4][17]  ( .D(n4420), .CLK(clk_in), .RSTB(n7114), .Q(
        \FIFO[4][17] ) );
  DFFARX1 \FIFO_reg[4][16]  ( .D(n4419), .CLK(clk_in), .RSTB(n7114), .Q(
        \FIFO[4][16] ) );
  DFFARX1 \FIFO_reg[4][15]  ( .D(n4418), .CLK(clk_in), .RSTB(n7114), .Q(
        \FIFO[4][15] ) );
  DFFARX1 \FIFO_reg[4][14]  ( .D(n4417), .CLK(clk_in), .RSTB(n7114), .Q(
        \FIFO[4][14] ) );
  DFFARX1 \FIFO_reg[4][13]  ( .D(n4416), .CLK(clk_in), .RSTB(n7114), .Q(
        \FIFO[4][13] ) );
  DFFARX1 \FIFO_reg[4][12]  ( .D(n4415), .CLK(clk_in), .RSTB(n7114), .Q(
        \FIFO[4][12] ) );
  DFFARX1 \FIFO_reg[4][11]  ( .D(n4414), .CLK(clk_in), .RSTB(n7114), .Q(
        \FIFO[4][11] ) );
  DFFARX1 \FIFO_reg[4][10]  ( .D(n4413), .CLK(clk_in), .RSTB(n7114), .Q(
        \FIFO[4][10] ) );
  DFFARX1 \FIFO_reg[4][9]  ( .D(n4412), .CLK(clk_in), .RSTB(n7115), .Q(
        \FIFO[4][9] ) );
  DFFARX1 \FIFO_reg[4][8]  ( .D(n4411), .CLK(clk_in), .RSTB(n7115), .Q(
        \FIFO[4][8] ) );
  DFFARX1 \FIFO_reg[4][7]  ( .D(n4410), .CLK(clk_in), .RSTB(n7115), .Q(
        \FIFO[4][7] ) );
  DFFARX1 \FIFO_reg[4][6]  ( .D(n4409), .CLK(clk_in), .RSTB(n7115), .Q(
        \FIFO[4][6] ) );
  DFFARX1 \FIFO_reg[4][5]  ( .D(n4408), .CLK(clk_in), .RSTB(n7115), .Q(
        \FIFO[4][5] ) );
  DFFARX1 \FIFO_reg[4][4]  ( .D(n4407), .CLK(clk_in), .RSTB(n7115), .Q(
        \FIFO[4][4] ) );
  DFFARX1 \FIFO_reg[4][3]  ( .D(n4406), .CLK(clk_in), .RSTB(n7115), .Q(
        \FIFO[4][3] ) );
  DFFARX1 \FIFO_reg[4][2]  ( .D(n4405), .CLK(clk_in), .RSTB(n7115), .Q(
        \FIFO[4][2] ) );
  DFFARX1 \FIFO_reg[4][1]  ( .D(n4404), .CLK(clk_in), .RSTB(n7115), .Q(
        \FIFO[4][1] ) );
  DFFARX1 \FIFO_reg[4][0]  ( .D(n4403), .CLK(clk_in), .RSTB(n7115), .Q(
        \FIFO[4][0] ) );
  DFFARX1 \FIFO_reg[5][31]  ( .D(n4402), .CLK(clk_in), .RSTB(n7115), .Q(
        \FIFO[5][31] ) );
  DFFARX1 \FIFO_reg[5][30]  ( .D(n4401), .CLK(clk_in), .RSTB(n7115), .Q(
        \FIFO[5][30] ) );
  DFFARX1 \FIFO_reg[5][29]  ( .D(n4400), .CLK(clk_in), .RSTB(n7115), .Q(
        \FIFO[5][29] ) );
  DFFARX1 \FIFO_reg[5][28]  ( .D(n4399), .CLK(clk_in), .RSTB(n7115), .Q(
        \FIFO[5][28] ) );
  DFFARX1 \FIFO_reg[5][27]  ( .D(n4398), .CLK(clk_in), .RSTB(n7115), .Q(
        \FIFO[5][27] ) );
  DFFARX1 \FIFO_reg[5][26]  ( .D(n4397), .CLK(clk_in), .RSTB(n7115), .Q(
        \FIFO[5][26] ) );
  DFFARX1 \FIFO_reg[5][25]  ( .D(n4396), .CLK(clk_in), .RSTB(n7115), .Q(
        \FIFO[5][25] ) );
  DFFARX1 \FIFO_reg[5][24]  ( .D(n4395), .CLK(clk_in), .RSTB(n7115), .Q(
        \FIFO[5][24] ) );
  DFFARX1 \FIFO_reg[5][23]  ( .D(n4394), .CLK(clk_in), .RSTB(n7116), .Q(
        \FIFO[5][23] ) );
  DFFARX1 \FIFO_reg[5][22]  ( .D(n4393), .CLK(clk_in), .RSTB(n7116), .Q(
        \FIFO[5][22] ) );
  DFFARX1 \FIFO_reg[5][21]  ( .D(n4392), .CLK(clk_in), .RSTB(n7116), .Q(
        \FIFO[5][21] ) );
  DFFARX1 \FIFO_reg[5][20]  ( .D(n4391), .CLK(clk_in), .RSTB(n7116), .Q(
        \FIFO[5][20] ) );
  DFFARX1 \FIFO_reg[5][19]  ( .D(n4390), .CLK(clk_in), .RSTB(n7116), .Q(
        \FIFO[5][19] ) );
  DFFARX1 \FIFO_reg[5][18]  ( .D(n4389), .CLK(clk_in), .RSTB(n7116), .Q(
        \FIFO[5][18] ) );
  DFFARX1 \FIFO_reg[5][17]  ( .D(n4388), .CLK(clk_in), .RSTB(n7116), .Q(
        \FIFO[5][17] ) );
  DFFARX1 \FIFO_reg[5][16]  ( .D(n4387), .CLK(clk_in), .RSTB(n7116), .Q(
        \FIFO[5][16] ) );
  DFFARX1 \FIFO_reg[5][15]  ( .D(n4386), .CLK(clk_in), .RSTB(n7116), .Q(
        \FIFO[5][15] ) );
  DFFARX1 \FIFO_reg[5][14]  ( .D(n4385), .CLK(clk_in), .RSTB(n7116), .Q(
        \FIFO[5][14] ) );
  DFFARX1 \FIFO_reg[5][13]  ( .D(n4384), .CLK(clk_in), .RSTB(n7116), .Q(
        \FIFO[5][13] ) );
  DFFARX1 \FIFO_reg[5][12]  ( .D(n4383), .CLK(clk_in), .RSTB(n7116), .Q(
        \FIFO[5][12] ) );
  DFFARX1 \FIFO_reg[5][11]  ( .D(n4382), .CLK(clk_in), .RSTB(n7116), .Q(
        \FIFO[5][11] ) );
  DFFARX1 \FIFO_reg[5][10]  ( .D(n4381), .CLK(clk_in), .RSTB(n7116), .Q(
        \FIFO[5][10] ) );
  DFFARX1 \FIFO_reg[5][9]  ( .D(n4380), .CLK(clk_in), .RSTB(n7116), .Q(
        \FIFO[5][9] ) );
  DFFARX1 \FIFO_reg[5][8]  ( .D(n4379), .CLK(clk_in), .RSTB(n7116), .Q(
        \FIFO[5][8] ) );
  DFFARX1 \FIFO_reg[5][7]  ( .D(n4378), .CLK(clk_in), .RSTB(n7116), .Q(
        \FIFO[5][7] ) );
  DFFARX1 \FIFO_reg[5][6]  ( .D(n4377), .CLK(clk_in), .RSTB(n7116), .Q(
        \FIFO[5][6] ) );
  DFFARX1 \FIFO_reg[5][5]  ( .D(n4376), .CLK(clk_in), .RSTB(n7117), .Q(
        \FIFO[5][5] ) );
  DFFARX1 \FIFO_reg[5][4]  ( .D(n4375), .CLK(clk_in), .RSTB(n7117), .Q(
        \FIFO[5][4] ) );
  DFFARX1 \FIFO_reg[5][3]  ( .D(n4374), .CLK(clk_in), .RSTB(n7117), .Q(
        \FIFO[5][3] ) );
  DFFARX1 \FIFO_reg[5][2]  ( .D(n4373), .CLK(clk_in), .RSTB(n7117), .Q(
        \FIFO[5][2] ) );
  DFFARX1 \FIFO_reg[5][1]  ( .D(n4372), .CLK(clk_in), .RSTB(n7117), .Q(
        \FIFO[5][1] ) );
  DFFARX1 \FIFO_reg[5][0]  ( .D(n4371), .CLK(clk_in), .RSTB(n7117), .Q(
        \FIFO[5][0] ) );
  DFFARX1 \FIFO_reg[6][31]  ( .D(n4370), .CLK(clk_in), .RSTB(n7117), .Q(
        \FIFO[6][31] ) );
  DFFARX1 \FIFO_reg[6][30]  ( .D(n4369), .CLK(clk_in), .RSTB(n7117), .Q(
        \FIFO[6][30] ) );
  DFFARX1 \FIFO_reg[6][29]  ( .D(n4368), .CLK(clk_in), .RSTB(n7117), .Q(
        \FIFO[6][29] ) );
  DFFARX1 \FIFO_reg[6][28]  ( .D(n4367), .CLK(clk_in), .RSTB(n7117), .Q(
        \FIFO[6][28] ) );
  DFFARX1 \FIFO_reg[6][27]  ( .D(n4366), .CLK(clk_in), .RSTB(n7117), .Q(
        \FIFO[6][27] ) );
  DFFARX1 \FIFO_reg[6][26]  ( .D(n4365), .CLK(clk_in), .RSTB(n7117), .Q(
        \FIFO[6][26] ) );
  DFFARX1 \FIFO_reg[6][25]  ( .D(n4364), .CLK(clk_in), .RSTB(n7117), .Q(
        \FIFO[6][25] ) );
  DFFARX1 \FIFO_reg[6][24]  ( .D(n4363), .CLK(clk_in), .RSTB(n7117), .Q(
        \FIFO[6][24] ) );
  DFFARX1 \FIFO_reg[6][23]  ( .D(n4362), .CLK(clk_in), .RSTB(n7117), .Q(
        \FIFO[6][23] ) );
  DFFARX1 \FIFO_reg[6][22]  ( .D(n4361), .CLK(clk_in), .RSTB(n7117), .Q(
        \FIFO[6][22] ) );
  DFFARX1 \FIFO_reg[6][21]  ( .D(n4360), .CLK(clk_in), .RSTB(n7117), .Q(
        \FIFO[6][21] ) );
  DFFARX1 \FIFO_reg[6][20]  ( .D(n4359), .CLK(clk_in), .RSTB(n7117), .Q(
        \FIFO[6][20] ) );
  DFFARX1 \FIFO_reg[6][19]  ( .D(n4358), .CLK(clk_in), .RSTB(n7118), .Q(
        \FIFO[6][19] ) );
  DFFARX1 \FIFO_reg[6][18]  ( .D(n4357), .CLK(clk_in), .RSTB(n7118), .Q(
        \FIFO[6][18] ) );
  DFFARX1 \FIFO_reg[6][17]  ( .D(n4356), .CLK(clk_in), .RSTB(n7118), .Q(
        \FIFO[6][17] ) );
  DFFARX1 \FIFO_reg[6][16]  ( .D(n4355), .CLK(clk_in), .RSTB(n7118), .Q(
        \FIFO[6][16] ) );
  DFFARX1 \FIFO_reg[6][15]  ( .D(n4354), .CLK(clk_in), .RSTB(n7118), .Q(
        \FIFO[6][15] ) );
  DFFARX1 \FIFO_reg[6][14]  ( .D(n4353), .CLK(clk_in), .RSTB(n7118), .Q(
        \FIFO[6][14] ) );
  DFFARX1 \FIFO_reg[6][13]  ( .D(n4352), .CLK(clk_in), .RSTB(n7118), .Q(
        \FIFO[6][13] ) );
  DFFARX1 \FIFO_reg[6][12]  ( .D(n4351), .CLK(clk_in), .RSTB(n7118), .Q(
        \FIFO[6][12] ) );
  DFFARX1 \FIFO_reg[6][11]  ( .D(n4350), .CLK(clk_in), .RSTB(n7118), .Q(
        \FIFO[6][11] ) );
  DFFARX1 \FIFO_reg[6][10]  ( .D(n4349), .CLK(clk_in), .RSTB(n7118), .Q(
        \FIFO[6][10] ) );
  DFFARX1 \FIFO_reg[6][9]  ( .D(n4348), .CLK(clk_in), .RSTB(n7118), .Q(
        \FIFO[6][9] ) );
  DFFARX1 \FIFO_reg[6][8]  ( .D(n4347), .CLK(clk_in), .RSTB(n7118), .Q(
        \FIFO[6][8] ) );
  DFFARX1 \FIFO_reg[6][7]  ( .D(n4346), .CLK(clk_in), .RSTB(n7118), .Q(
        \FIFO[6][7] ) );
  DFFARX1 \FIFO_reg[6][6]  ( .D(n4345), .CLK(clk_in), .RSTB(n7118), .Q(
        \FIFO[6][6] ) );
  DFFARX1 \FIFO_reg[6][5]  ( .D(n4344), .CLK(clk_in), .RSTB(n7118), .Q(
        \FIFO[6][5] ) );
  DFFARX1 \FIFO_reg[6][4]  ( .D(n4343), .CLK(clk_in), .RSTB(n7118), .Q(
        \FIFO[6][4] ) );
  DFFARX1 \FIFO_reg[6][3]  ( .D(n4342), .CLK(clk_in), .RSTB(n7118), .Q(
        \FIFO[6][3] ) );
  DFFARX1 \FIFO_reg[6][2]  ( .D(n4341), .CLK(clk_in), .RSTB(n7118), .Q(
        \FIFO[6][2] ) );
  DFFARX1 \FIFO_reg[6][1]  ( .D(n4340), .CLK(clk_in), .RSTB(n7119), .Q(
        \FIFO[6][1] ) );
  DFFARX1 \FIFO_reg[6][0]  ( .D(n4339), .CLK(clk_in), .RSTB(n7119), .Q(
        \FIFO[6][0] ) );
  DFFARX1 \FIFO_reg[7][31]  ( .D(n4338), .CLK(clk_in), .RSTB(n7119), .Q(
        \FIFO[7][31] ) );
  DFFARX1 \FIFO_reg[7][30]  ( .D(n4337), .CLK(clk_in), .RSTB(n7119), .Q(
        \FIFO[7][30] ) );
  DFFARX1 \FIFO_reg[7][29]  ( .D(n4336), .CLK(clk_in), .RSTB(n7119), .Q(
        \FIFO[7][29] ) );
  DFFARX1 \FIFO_reg[7][28]  ( .D(n4335), .CLK(clk_in), .RSTB(n7119), .Q(
        \FIFO[7][28] ) );
  DFFARX1 \FIFO_reg[7][27]  ( .D(n4334), .CLK(clk_in), .RSTB(n7119), .Q(
        \FIFO[7][27] ) );
  DFFARX1 \FIFO_reg[7][26]  ( .D(n4333), .CLK(clk_in), .RSTB(n7119), .Q(
        \FIFO[7][26] ) );
  DFFARX1 \FIFO_reg[7][25]  ( .D(n4332), .CLK(clk_in), .RSTB(n7119), .Q(
        \FIFO[7][25] ) );
  DFFARX1 \FIFO_reg[7][24]  ( .D(n4331), .CLK(clk_in), .RSTB(n7119), .Q(
        \FIFO[7][24] ) );
  DFFARX1 \FIFO_reg[7][23]  ( .D(n4330), .CLK(clk_in), .RSTB(n7119), .Q(
        \FIFO[7][23] ) );
  DFFARX1 \FIFO_reg[7][22]  ( .D(n4329), .CLK(clk_in), .RSTB(n7119), .Q(
        \FIFO[7][22] ) );
  DFFARX1 \FIFO_reg[7][21]  ( .D(n4328), .CLK(clk_in), .RSTB(n7119), .Q(
        \FIFO[7][21] ) );
  DFFARX1 \FIFO_reg[7][20]  ( .D(n4327), .CLK(clk_in), .RSTB(n7119), .Q(
        \FIFO[7][20] ) );
  DFFARX1 \FIFO_reg[7][19]  ( .D(n4326), .CLK(clk_in), .RSTB(n7119), .Q(
        \FIFO[7][19] ) );
  DFFARX1 \FIFO_reg[7][18]  ( .D(n4325), .CLK(clk_in), .RSTB(n7119), .Q(
        \FIFO[7][18] ) );
  DFFARX1 \FIFO_reg[7][17]  ( .D(n4324), .CLK(clk_in), .RSTB(n7119), .Q(
        \FIFO[7][17] ) );
  DFFARX1 \FIFO_reg[7][16]  ( .D(n4323), .CLK(clk_in), .RSTB(n7119), .Q(
        \FIFO[7][16] ) );
  DFFARX1 \FIFO_reg[7][15]  ( .D(n4322), .CLK(clk_in), .RSTB(n7120), .Q(
        \FIFO[7][15] ) );
  DFFARX1 \FIFO_reg[7][14]  ( .D(n4321), .CLK(clk_in), .RSTB(n7120), .Q(
        \FIFO[7][14] ) );
  DFFARX1 \FIFO_reg[7][13]  ( .D(n4320), .CLK(clk_in), .RSTB(n7120), .Q(
        \FIFO[7][13] ) );
  DFFARX1 \FIFO_reg[7][12]  ( .D(n4319), .CLK(clk_in), .RSTB(n7120), .Q(
        \FIFO[7][12] ) );
  DFFARX1 \FIFO_reg[7][11]  ( .D(n4318), .CLK(clk_in), .RSTB(n7120), .Q(
        \FIFO[7][11] ) );
  DFFARX1 \FIFO_reg[7][10]  ( .D(n4317), .CLK(clk_in), .RSTB(n7120), .Q(
        \FIFO[7][10] ) );
  DFFARX1 \FIFO_reg[7][9]  ( .D(n4316), .CLK(clk_in), .RSTB(n7120), .Q(
        \FIFO[7][9] ) );
  DFFARX1 \FIFO_reg[7][8]  ( .D(n4315), .CLK(clk_in), .RSTB(n7120), .Q(
        \FIFO[7][8] ) );
  DFFARX1 \FIFO_reg[7][7]  ( .D(n4314), .CLK(clk_in), .RSTB(n7120), .Q(
        \FIFO[7][7] ) );
  DFFARX1 \FIFO_reg[7][6]  ( .D(n4313), .CLK(clk_in), .RSTB(n7120), .Q(
        \FIFO[7][6] ) );
  DFFARX1 \FIFO_reg[7][5]  ( .D(n4312), .CLK(clk_in), .RSTB(n7120), .Q(
        \FIFO[7][5] ) );
  DFFARX1 \FIFO_reg[7][4]  ( .D(n4311), .CLK(clk_in), .RSTB(n7120), .Q(
        \FIFO[7][4] ) );
  DFFARX1 \FIFO_reg[7][3]  ( .D(n4310), .CLK(clk_in), .RSTB(n7120), .Q(
        \FIFO[7][3] ) );
  DFFARX1 \FIFO_reg[7][2]  ( .D(n4309), .CLK(clk_in), .RSTB(n7120), .Q(
        \FIFO[7][2] ) );
  DFFARX1 \FIFO_reg[7][1]  ( .D(n4308), .CLK(clk_in), .RSTB(n7120), .Q(
        \FIFO[7][1] ) );
  DFFARX1 \FIFO_reg[7][0]  ( .D(n4307), .CLK(clk_in), .RSTB(n7120), .Q(
        \FIFO[7][0] ) );
  DFFARX1 \FIFO_reg[8][31]  ( .D(n4306), .CLK(clk_in), .RSTB(n7120), .Q(
        \FIFO[8][31] ) );
  DFFARX1 \FIFO_reg[8][30]  ( .D(n4305), .CLK(clk_in), .RSTB(n7120), .Q(
        \FIFO[8][30] ) );
  DFFARX1 \FIFO_reg[8][29]  ( .D(n4304), .CLK(clk_in), .RSTB(n7121), .Q(
        \FIFO[8][29] ) );
  DFFARX1 \FIFO_reg[8][28]  ( .D(n4303), .CLK(clk_in), .RSTB(n7121), .Q(
        \FIFO[8][28] ) );
  DFFARX1 \FIFO_reg[8][27]  ( .D(n4302), .CLK(clk_in), .RSTB(n7121), .Q(
        \FIFO[8][27] ) );
  DFFARX1 \FIFO_reg[8][26]  ( .D(n4301), .CLK(clk_in), .RSTB(n7121), .Q(
        \FIFO[8][26] ) );
  DFFARX1 \FIFO_reg[8][25]  ( .D(n4300), .CLK(clk_in), .RSTB(n7121), .Q(
        \FIFO[8][25] ) );
  DFFARX1 \FIFO_reg[8][24]  ( .D(n4299), .CLK(clk_in), .RSTB(n7121), .Q(
        \FIFO[8][24] ) );
  DFFARX1 \FIFO_reg[8][23]  ( .D(n4298), .CLK(clk_in), .RSTB(n7121), .Q(
        \FIFO[8][23] ) );
  DFFARX1 \FIFO_reg[8][22]  ( .D(n4297), .CLK(clk_in), .RSTB(n7121), .Q(
        \FIFO[8][22] ) );
  DFFARX1 \FIFO_reg[8][21]  ( .D(n4296), .CLK(clk_in), .RSTB(n7121), .Q(
        \FIFO[8][21] ) );
  DFFARX1 \FIFO_reg[8][20]  ( .D(n4295), .CLK(clk_in), .RSTB(n7121), .Q(
        \FIFO[8][20] ) );
  DFFARX1 \FIFO_reg[8][19]  ( .D(n4294), .CLK(clk_in), .RSTB(n7121), .Q(
        \FIFO[8][19] ) );
  DFFARX1 \FIFO_reg[8][18]  ( .D(n4293), .CLK(clk_in), .RSTB(n7121), .Q(
        \FIFO[8][18] ) );
  DFFARX1 \FIFO_reg[8][17]  ( .D(n4292), .CLK(clk_in), .RSTB(n7121), .Q(
        \FIFO[8][17] ) );
  DFFARX1 \FIFO_reg[8][16]  ( .D(n4291), .CLK(clk_in), .RSTB(n7121), .Q(
        \FIFO[8][16] ) );
  DFFARX1 \FIFO_reg[8][15]  ( .D(n4290), .CLK(clk_in), .RSTB(n7121), .Q(
        \FIFO[8][15] ) );
  DFFARX1 \FIFO_reg[8][14]  ( .D(n4289), .CLK(clk_in), .RSTB(n7121), .Q(
        \FIFO[8][14] ) );
  DFFARX1 \FIFO_reg[8][13]  ( .D(n4288), .CLK(clk_in), .RSTB(n7121), .Q(
        \FIFO[8][13] ) );
  DFFARX1 \FIFO_reg[8][12]  ( .D(n4287), .CLK(clk_in), .RSTB(n7121), .Q(
        \FIFO[8][12] ) );
  DFFARX1 \FIFO_reg[8][11]  ( .D(n4286), .CLK(clk_in), .RSTB(n7122), .Q(
        \FIFO[8][11] ) );
  DFFARX1 \FIFO_reg[8][10]  ( .D(n4285), .CLK(clk_in), .RSTB(n7122), .Q(
        \FIFO[8][10] ) );
  DFFARX1 \FIFO_reg[8][9]  ( .D(n4284), .CLK(clk_in), .RSTB(n7122), .Q(
        \FIFO[8][9] ) );
  DFFARX1 \FIFO_reg[8][8]  ( .D(n4283), .CLK(clk_in), .RSTB(n7122), .Q(
        \FIFO[8][8] ) );
  DFFARX1 \FIFO_reg[8][7]  ( .D(n4282), .CLK(clk_in), .RSTB(n7122), .Q(
        \FIFO[8][7] ) );
  DFFARX1 \FIFO_reg[8][6]  ( .D(n4281), .CLK(clk_in), .RSTB(n7122), .Q(
        \FIFO[8][6] ) );
  DFFARX1 \FIFO_reg[8][5]  ( .D(n4280), .CLK(clk_in), .RSTB(n7122), .Q(
        \FIFO[8][5] ) );
  DFFARX1 \FIFO_reg[8][4]  ( .D(n4279), .CLK(clk_in), .RSTB(n7122), .Q(
        \FIFO[8][4] ) );
  DFFARX1 \FIFO_reg[8][3]  ( .D(n4278), .CLK(clk_in), .RSTB(n7122), .Q(
        \FIFO[8][3] ) );
  DFFARX1 \FIFO_reg[8][2]  ( .D(n4277), .CLK(clk_in), .RSTB(n7122), .Q(
        \FIFO[8][2] ) );
  DFFARX1 \FIFO_reg[8][1]  ( .D(n4276), .CLK(clk_in), .RSTB(n7122), .Q(
        \FIFO[8][1] ) );
  DFFARX1 \FIFO_reg[8][0]  ( .D(n4275), .CLK(clk_in), .RSTB(n7122), .Q(
        \FIFO[8][0] ) );
  DFFARX1 \FIFO_reg[9][31]  ( .D(n4274), .CLK(clk_in), .RSTB(n7122), .Q(
        \FIFO[9][31] ) );
  DFFARX1 \FIFO_reg[9][30]  ( .D(n4273), .CLK(clk_in), .RSTB(n7122), .Q(
        \FIFO[9][30] ) );
  DFFARX1 \FIFO_reg[9][29]  ( .D(n4272), .CLK(clk_in), .RSTB(n7122), .Q(
        \FIFO[9][29] ) );
  DFFARX1 \FIFO_reg[9][28]  ( .D(n4271), .CLK(clk_in), .RSTB(n7122), .Q(
        \FIFO[9][28] ) );
  DFFARX1 \FIFO_reg[9][27]  ( .D(n4270), .CLK(clk_in), .RSTB(n7122), .Q(
        \FIFO[9][27] ) );
  DFFARX1 \FIFO_reg[9][26]  ( .D(n4269), .CLK(clk_in), .RSTB(n7122), .Q(
        \FIFO[9][26] ) );
  DFFARX1 \FIFO_reg[9][25]  ( .D(n4268), .CLK(clk_in), .RSTB(n7123), .Q(
        \FIFO[9][25] ) );
  DFFARX1 \FIFO_reg[9][24]  ( .D(n4267), .CLK(clk_in), .RSTB(n7123), .Q(
        \FIFO[9][24] ) );
  DFFARX1 \FIFO_reg[9][23]  ( .D(n4266), .CLK(clk_in), .RSTB(n7123), .Q(
        \FIFO[9][23] ) );
  DFFARX1 \FIFO_reg[9][22]  ( .D(n4265), .CLK(clk_in), .RSTB(n7123), .Q(
        \FIFO[9][22] ) );
  DFFARX1 \FIFO_reg[9][21]  ( .D(n4264), .CLK(clk_in), .RSTB(n7123), .Q(
        \FIFO[9][21] ) );
  DFFARX1 \FIFO_reg[9][20]  ( .D(n4263), .CLK(clk_in), .RSTB(n7123), .Q(
        \FIFO[9][20] ) );
  DFFARX1 \FIFO_reg[9][19]  ( .D(n4262), .CLK(clk_in), .RSTB(n7123), .Q(
        \FIFO[9][19] ) );
  DFFARX1 \FIFO_reg[9][18]  ( .D(n4261), .CLK(clk_in), .RSTB(n7123), .Q(
        \FIFO[9][18] ) );
  DFFARX1 \FIFO_reg[9][17]  ( .D(n4260), .CLK(clk_in), .RSTB(n7123), .Q(
        \FIFO[9][17] ) );
  DFFARX1 \FIFO_reg[9][16]  ( .D(n4259), .CLK(clk_in), .RSTB(n7123), .Q(
        \FIFO[9][16] ) );
  DFFARX1 \FIFO_reg[9][15]  ( .D(n4258), .CLK(clk_in), .RSTB(n7123), .Q(
        \FIFO[9][15] ) );
  DFFARX1 \FIFO_reg[9][14]  ( .D(n4257), .CLK(clk_in), .RSTB(n7123), .Q(
        \FIFO[9][14] ) );
  DFFARX1 \FIFO_reg[9][13]  ( .D(n4256), .CLK(clk_in), .RSTB(n7123), .Q(
        \FIFO[9][13] ) );
  DFFARX1 \FIFO_reg[9][12]  ( .D(n4255), .CLK(clk_in), .RSTB(n7123), .Q(
        \FIFO[9][12] ) );
  DFFARX1 \FIFO_reg[9][11]  ( .D(n4254), .CLK(clk_in), .RSTB(n7123), .Q(
        \FIFO[9][11] ) );
  DFFARX1 \FIFO_reg[9][10]  ( .D(n4253), .CLK(clk_in), .RSTB(n7123), .Q(
        \FIFO[9][10] ) );
  DFFARX1 \FIFO_reg[9][9]  ( .D(n4252), .CLK(clk_in), .RSTB(n7123), .Q(
        \FIFO[9][9] ) );
  DFFARX1 \FIFO_reg[9][8]  ( .D(n4251), .CLK(clk_in), .RSTB(n7123), .Q(
        \FIFO[9][8] ) );
  DFFARX1 \FIFO_reg[9][7]  ( .D(n4250), .CLK(clk_in), .RSTB(n7124), .Q(
        \FIFO[9][7] ) );
  DFFARX1 \FIFO_reg[9][6]  ( .D(n4249), .CLK(clk_in), .RSTB(n7124), .Q(
        \FIFO[9][6] ) );
  DFFARX1 \FIFO_reg[9][5]  ( .D(n4248), .CLK(clk_in), .RSTB(n7124), .Q(
        \FIFO[9][5] ) );
  DFFARX1 \FIFO_reg[9][4]  ( .D(n4247), .CLK(clk_in), .RSTB(n7124), .Q(
        \FIFO[9][4] ) );
  DFFARX1 \FIFO_reg[9][3]  ( .D(n4246), .CLK(clk_in), .RSTB(n7124), .Q(
        \FIFO[9][3] ) );
  DFFARX1 \FIFO_reg[9][2]  ( .D(n4245), .CLK(clk_in), .RSTB(n7124), .Q(
        \FIFO[9][2] ) );
  DFFARX1 \FIFO_reg[9][1]  ( .D(n4244), .CLK(clk_in), .RSTB(n7124), .Q(
        \FIFO[9][1] ) );
  DFFARX1 \FIFO_reg[9][0]  ( .D(n4243), .CLK(clk_in), .RSTB(n7124), .Q(
        \FIFO[9][0] ) );
  DFFARX1 \FIFO_reg[10][31]  ( .D(n4242), .CLK(clk_in), .RSTB(n7124), .Q(
        \FIFO[10][31] ) );
  DFFARX1 \FIFO_reg[10][30]  ( .D(n4241), .CLK(clk_in), .RSTB(n7124), .Q(
        \FIFO[10][30] ) );
  DFFARX1 \FIFO_reg[10][29]  ( .D(n4240), .CLK(clk_in), .RSTB(n7124), .Q(
        \FIFO[10][29] ) );
  DFFARX1 \FIFO_reg[10][28]  ( .D(n4239), .CLK(clk_in), .RSTB(n7124), .Q(
        \FIFO[10][28] ) );
  DFFARX1 \FIFO_reg[10][27]  ( .D(n4238), .CLK(clk_in), .RSTB(n7124), .Q(
        \FIFO[10][27] ) );
  DFFARX1 \FIFO_reg[10][26]  ( .D(n4237), .CLK(clk_in), .RSTB(n7124), .Q(
        \FIFO[10][26] ) );
  DFFARX1 \FIFO_reg[10][25]  ( .D(n4236), .CLK(clk_in), .RSTB(n7124), .Q(
        \FIFO[10][25] ) );
  DFFARX1 \FIFO_reg[10][24]  ( .D(n4235), .CLK(clk_in), .RSTB(n7124), .Q(
        \FIFO[10][24] ) );
  DFFARX1 \FIFO_reg[10][23]  ( .D(n4234), .CLK(clk_in), .RSTB(n7124), .Q(
        \FIFO[10][23] ) );
  DFFARX1 \FIFO_reg[10][22]  ( .D(n4233), .CLK(clk_in), .RSTB(n7124), .Q(
        \FIFO[10][22] ) );
  DFFARX1 \FIFO_reg[10][21]  ( .D(n4232), .CLK(clk_in), .RSTB(n7125), .Q(
        \FIFO[10][21] ) );
  DFFARX1 \FIFO_reg[10][20]  ( .D(n4231), .CLK(clk_in), .RSTB(n7125), .Q(
        \FIFO[10][20] ) );
  DFFARX1 \FIFO_reg[10][19]  ( .D(n4230), .CLK(clk_in), .RSTB(n7125), .Q(
        \FIFO[10][19] ) );
  DFFARX1 \FIFO_reg[10][18]  ( .D(n4229), .CLK(clk_in), .RSTB(n7125), .Q(
        \FIFO[10][18] ) );
  DFFARX1 \FIFO_reg[10][17]  ( .D(n4228), .CLK(clk_in), .RSTB(n7125), .Q(
        \FIFO[10][17] ) );
  DFFARX1 \FIFO_reg[10][16]  ( .D(n4227), .CLK(clk_in), .RSTB(n7125), .Q(
        \FIFO[10][16] ) );
  DFFARX1 \FIFO_reg[10][15]  ( .D(n4226), .CLK(clk_in), .RSTB(n7125), .Q(
        \FIFO[10][15] ) );
  DFFARX1 \FIFO_reg[10][14]  ( .D(n4225), .CLK(clk_in), .RSTB(n7125), .Q(
        \FIFO[10][14] ) );
  DFFARX1 \FIFO_reg[10][13]  ( .D(n4224), .CLK(clk_in), .RSTB(n7125), .Q(
        \FIFO[10][13] ) );
  DFFARX1 \FIFO_reg[10][12]  ( .D(n4223), .CLK(clk_in), .RSTB(n7125), .Q(
        \FIFO[10][12] ) );
  DFFARX1 \FIFO_reg[10][11]  ( .D(n4222), .CLK(clk_in), .RSTB(n7125), .Q(
        \FIFO[10][11] ) );
  DFFARX1 \FIFO_reg[10][10]  ( .D(n4221), .CLK(clk_in), .RSTB(n7125), .Q(
        \FIFO[10][10] ) );
  DFFARX1 \FIFO_reg[10][9]  ( .D(n4220), .CLK(clk_in), .RSTB(n7125), .Q(
        \FIFO[10][9] ) );
  DFFARX1 \FIFO_reg[10][8]  ( .D(n4219), .CLK(clk_in), .RSTB(n7125), .Q(
        \FIFO[10][8] ) );
  DFFARX1 \FIFO_reg[10][7]  ( .D(n4218), .CLK(clk_in), .RSTB(n7125), .Q(
        \FIFO[10][7] ) );
  DFFARX1 \FIFO_reg[10][6]  ( .D(n4217), .CLK(clk_in), .RSTB(n7125), .Q(
        \FIFO[10][6] ) );
  DFFARX1 \FIFO_reg[10][5]  ( .D(n4216), .CLK(clk_in), .RSTB(n7125), .Q(
        \FIFO[10][5] ) );
  DFFARX1 \FIFO_reg[10][4]  ( .D(n4215), .CLK(clk_in), .RSTB(n7125), .Q(
        \FIFO[10][4] ) );
  DFFARX1 \FIFO_reg[10][3]  ( .D(n4214), .CLK(clk_in), .RSTB(n7126), .Q(
        \FIFO[10][3] ) );
  DFFARX1 \FIFO_reg[10][2]  ( .D(n4213), .CLK(clk_in), .RSTB(n7126), .Q(
        \FIFO[10][2] ) );
  DFFARX1 \FIFO_reg[10][1]  ( .D(n4212), .CLK(clk_in), .RSTB(n7126), .Q(
        \FIFO[10][1] ) );
  DFFARX1 \FIFO_reg[10][0]  ( .D(n4211), .CLK(clk_in), .RSTB(n7126), .Q(
        \FIFO[10][0] ) );
  DFFARX1 \FIFO_reg[11][31]  ( .D(n4210), .CLK(clk_in), .RSTB(n7126), .Q(
        \FIFO[11][31] ) );
  DFFARX1 \FIFO_reg[11][30]  ( .D(n4209), .CLK(clk_in), .RSTB(n7126), .Q(
        \FIFO[11][30] ) );
  DFFARX1 \FIFO_reg[11][29]  ( .D(n4208), .CLK(clk_in), .RSTB(n7126), .Q(
        \FIFO[11][29] ) );
  DFFARX1 \FIFO_reg[11][28]  ( .D(n4207), .CLK(clk_in), .RSTB(n7126), .Q(
        \FIFO[11][28] ) );
  DFFARX1 \FIFO_reg[11][27]  ( .D(n4206), .CLK(clk_in), .RSTB(n7126), .Q(
        \FIFO[11][27] ) );
  DFFARX1 \FIFO_reg[11][26]  ( .D(n4205), .CLK(clk_in), .RSTB(n7126), .Q(
        \FIFO[11][26] ) );
  DFFARX1 \FIFO_reg[11][25]  ( .D(n4204), .CLK(clk_in), .RSTB(n7126), .Q(
        \FIFO[11][25] ) );
  DFFARX1 \FIFO_reg[11][24]  ( .D(n4203), .CLK(clk_in), .RSTB(n7126), .Q(
        \FIFO[11][24] ) );
  DFFARX1 \FIFO_reg[11][23]  ( .D(n4202), .CLK(clk_in), .RSTB(n7126), .Q(
        \FIFO[11][23] ) );
  DFFARX1 \FIFO_reg[11][22]  ( .D(n4201), .CLK(clk_in), .RSTB(n7126), .Q(
        \FIFO[11][22] ) );
  DFFARX1 \FIFO_reg[11][21]  ( .D(n4200), .CLK(clk_in), .RSTB(n7126), .Q(
        \FIFO[11][21] ) );
  DFFARX1 \FIFO_reg[11][20]  ( .D(n4199), .CLK(clk_in), .RSTB(n7126), .Q(
        \FIFO[11][20] ) );
  DFFARX1 \FIFO_reg[11][19]  ( .D(n4198), .CLK(clk_in), .RSTB(n7126), .Q(
        \FIFO[11][19] ) );
  DFFARX1 \FIFO_reg[11][18]  ( .D(n4197), .CLK(clk_in), .RSTB(n7126), .Q(
        \FIFO[11][18] ) );
  DFFARX1 \FIFO_reg[11][17]  ( .D(n4196), .CLK(clk_in), .RSTB(n7127), .Q(
        \FIFO[11][17] ) );
  DFFARX1 \FIFO_reg[11][16]  ( .D(n4195), .CLK(clk_in), .RSTB(n7127), .Q(
        \FIFO[11][16] ) );
  DFFARX1 \FIFO_reg[11][15]  ( .D(n4194), .CLK(clk_in), .RSTB(n7127), .Q(
        \FIFO[11][15] ) );
  DFFARX1 \FIFO_reg[11][14]  ( .D(n4193), .CLK(clk_in), .RSTB(n7127), .Q(
        \FIFO[11][14] ) );
  DFFARX1 \FIFO_reg[11][13]  ( .D(n4192), .CLK(clk_in), .RSTB(n7127), .Q(
        \FIFO[11][13] ) );
  DFFARX1 \FIFO_reg[11][12]  ( .D(n4191), .CLK(clk_in), .RSTB(n7127), .Q(
        \FIFO[11][12] ) );
  DFFARX1 \FIFO_reg[11][11]  ( .D(n4190), .CLK(clk_in), .RSTB(n7127), .Q(
        \FIFO[11][11] ) );
  DFFARX1 \FIFO_reg[11][10]  ( .D(n4189), .CLK(clk_in), .RSTB(n7127), .Q(
        \FIFO[11][10] ) );
  DFFARX1 \FIFO_reg[11][9]  ( .D(n4188), .CLK(clk_in), .RSTB(n7127), .Q(
        \FIFO[11][9] ) );
  DFFARX1 \FIFO_reg[11][8]  ( .D(n4187), .CLK(clk_in), .RSTB(n7127), .Q(
        \FIFO[11][8] ) );
  DFFARX1 \FIFO_reg[11][7]  ( .D(n4186), .CLK(clk_in), .RSTB(n7127), .Q(
        \FIFO[11][7] ) );
  DFFARX1 \FIFO_reg[11][6]  ( .D(n4185), .CLK(clk_in), .RSTB(n7127), .Q(
        \FIFO[11][6] ) );
  DFFARX1 \FIFO_reg[11][5]  ( .D(n4184), .CLK(clk_in), .RSTB(n7127), .Q(
        \FIFO[11][5] ) );
  DFFARX1 \FIFO_reg[11][4]  ( .D(n4183), .CLK(clk_in), .RSTB(n7127), .Q(
        \FIFO[11][4] ) );
  DFFARX1 \FIFO_reg[11][3]  ( .D(n4182), .CLK(clk_in), .RSTB(n7127), .Q(
        \FIFO[11][3] ) );
  DFFARX1 \FIFO_reg[11][2]  ( .D(n4181), .CLK(clk_in), .RSTB(n7127), .Q(
        \FIFO[11][2] ) );
  DFFARX1 \FIFO_reg[11][1]  ( .D(n4180), .CLK(clk_in), .RSTB(n7127), .Q(
        \FIFO[11][1] ) );
  DFFARX1 \FIFO_reg[11][0]  ( .D(n4179), .CLK(clk_in), .RSTB(n7127), .Q(
        \FIFO[11][0] ) );
  DFFARX1 \FIFO_reg[12][31]  ( .D(n4178), .CLK(clk_in), .RSTB(n7128), .Q(
        \FIFO[12][31] ) );
  DFFARX1 \FIFO_reg[12][30]  ( .D(n4177), .CLK(clk_in), .RSTB(n7128), .Q(
        \FIFO[12][30] ) );
  DFFARX1 \FIFO_reg[12][29]  ( .D(n4176), .CLK(clk_in), .RSTB(n7128), .Q(
        \FIFO[12][29] ) );
  DFFARX1 \FIFO_reg[12][28]  ( .D(n4175), .CLK(clk_in), .RSTB(n7128), .Q(
        \FIFO[12][28] ) );
  DFFARX1 \FIFO_reg[12][27]  ( .D(n4174), .CLK(clk_in), .RSTB(n7128), .Q(
        \FIFO[12][27] ) );
  DFFARX1 \FIFO_reg[12][26]  ( .D(n4173), .CLK(clk_in), .RSTB(n7128), .Q(
        \FIFO[12][26] ) );
  DFFARX1 \FIFO_reg[12][25]  ( .D(n4172), .CLK(clk_in), .RSTB(n7128), .Q(
        \FIFO[12][25] ) );
  DFFARX1 \FIFO_reg[12][24]  ( .D(n4171), .CLK(clk_in), .RSTB(n7128), .Q(
        \FIFO[12][24] ) );
  DFFARX1 \FIFO_reg[12][23]  ( .D(n4170), .CLK(clk_in), .RSTB(n7128), .Q(
        \FIFO[12][23] ) );
  DFFARX1 \FIFO_reg[12][22]  ( .D(n4169), .CLK(clk_in), .RSTB(n7128), .Q(
        \FIFO[12][22] ) );
  DFFARX1 \FIFO_reg[12][21]  ( .D(n4168), .CLK(clk_in), .RSTB(n7128), .Q(
        \FIFO[12][21] ) );
  DFFARX1 \FIFO_reg[12][20]  ( .D(n4167), .CLK(clk_in), .RSTB(n7128), .Q(
        \FIFO[12][20] ) );
  DFFARX1 \FIFO_reg[12][19]  ( .D(n4166), .CLK(clk_in), .RSTB(n7128), .Q(
        \FIFO[12][19] ) );
  DFFARX1 \FIFO_reg[12][18]  ( .D(n4165), .CLK(clk_in), .RSTB(n7128), .Q(
        \FIFO[12][18] ) );
  DFFARX1 \FIFO_reg[12][17]  ( .D(n4164), .CLK(clk_in), .RSTB(n7128), .Q(
        \FIFO[12][17] ) );
  DFFARX1 \FIFO_reg[12][16]  ( .D(n4163), .CLK(clk_in), .RSTB(n7128), .Q(
        \FIFO[12][16] ) );
  DFFARX1 \FIFO_reg[12][15]  ( .D(n4162), .CLK(clk_in), .RSTB(n7128), .Q(
        \FIFO[12][15] ) );
  DFFARX1 \FIFO_reg[12][14]  ( .D(n4161), .CLK(clk_in), .RSTB(n7128), .Q(
        \FIFO[12][14] ) );
  DFFARX1 \FIFO_reg[12][13]  ( .D(n4160), .CLK(clk_in), .RSTB(n7129), .Q(
        \FIFO[12][13] ) );
  DFFARX1 \FIFO_reg[12][12]  ( .D(n4159), .CLK(clk_in), .RSTB(n7129), .Q(
        \FIFO[12][12] ) );
  DFFARX1 \FIFO_reg[12][11]  ( .D(n4158), .CLK(clk_in), .RSTB(n7129), .Q(
        \FIFO[12][11] ) );
  DFFARX1 \FIFO_reg[12][10]  ( .D(n4157), .CLK(clk_in), .RSTB(n7129), .Q(
        \FIFO[12][10] ) );
  DFFARX1 \FIFO_reg[12][9]  ( .D(n4156), .CLK(clk_in), .RSTB(n7129), .Q(
        \FIFO[12][9] ) );
  DFFARX1 \FIFO_reg[12][8]  ( .D(n4155), .CLK(clk_in), .RSTB(n7129), .Q(
        \FIFO[12][8] ) );
  DFFARX1 \FIFO_reg[12][7]  ( .D(n4154), .CLK(clk_in), .RSTB(n7129), .Q(
        \FIFO[12][7] ) );
  DFFARX1 \FIFO_reg[12][6]  ( .D(n4153), .CLK(clk_in), .RSTB(n7129), .Q(
        \FIFO[12][6] ) );
  DFFARX1 \FIFO_reg[12][5]  ( .D(n4152), .CLK(clk_in), .RSTB(n7129), .Q(
        \FIFO[12][5] ) );
  DFFARX1 \FIFO_reg[12][4]  ( .D(n4151), .CLK(clk_in), .RSTB(n7129), .Q(
        \FIFO[12][4] ) );
  DFFARX1 \FIFO_reg[12][3]  ( .D(n4150), .CLK(clk_in), .RSTB(n7129), .Q(
        \FIFO[12][3] ) );
  DFFARX1 \FIFO_reg[12][2]  ( .D(n4149), .CLK(clk_in), .RSTB(n7129), .Q(
        \FIFO[12][2] ) );
  DFFARX1 \FIFO_reg[12][1]  ( .D(n4148), .CLK(clk_in), .RSTB(n7129), .Q(
        \FIFO[12][1] ) );
  DFFARX1 \FIFO_reg[12][0]  ( .D(n4147), .CLK(clk_in), .RSTB(n7129), .Q(
        \FIFO[12][0] ) );
  DFFARX1 \FIFO_reg[13][31]  ( .D(n4146), .CLK(clk_in), .RSTB(n7129), .Q(
        \FIFO[13][31] ) );
  DFFARX1 \FIFO_reg[13][30]  ( .D(n4145), .CLK(clk_in), .RSTB(n7129), .Q(
        \FIFO[13][30] ) );
  DFFARX1 \FIFO_reg[13][29]  ( .D(n4144), .CLK(clk_in), .RSTB(n7129), .Q(
        \FIFO[13][29] ) );
  DFFARX1 \FIFO_reg[13][28]  ( .D(n4143), .CLK(clk_in), .RSTB(n7129), .Q(
        \FIFO[13][28] ) );
  DFFARX1 \FIFO_reg[13][27]  ( .D(n4142), .CLK(clk_in), .RSTB(n7130), .Q(
        \FIFO[13][27] ) );
  DFFARX1 \FIFO_reg[13][26]  ( .D(n4141), .CLK(clk_in), .RSTB(n7130), .Q(
        \FIFO[13][26] ) );
  DFFARX1 \FIFO_reg[13][25]  ( .D(n4140), .CLK(clk_in), .RSTB(n7130), .Q(
        \FIFO[13][25] ) );
  DFFARX1 \FIFO_reg[13][24]  ( .D(n4139), .CLK(clk_in), .RSTB(n7130), .Q(
        \FIFO[13][24] ) );
  DFFARX1 \FIFO_reg[13][23]  ( .D(n4138), .CLK(clk_in), .RSTB(n7130), .Q(
        \FIFO[13][23] ) );
  DFFARX1 \FIFO_reg[13][22]  ( .D(n4137), .CLK(clk_in), .RSTB(n7130), .Q(
        \FIFO[13][22] ) );
  DFFARX1 \FIFO_reg[13][21]  ( .D(n4136), .CLK(clk_in), .RSTB(n7130), .Q(
        \FIFO[13][21] ) );
  DFFARX1 \FIFO_reg[13][20]  ( .D(n4135), .CLK(clk_in), .RSTB(n7130), .Q(
        \FIFO[13][20] ) );
  DFFARX1 \FIFO_reg[13][19]  ( .D(n4134), .CLK(clk_in), .RSTB(n7130), .Q(
        \FIFO[13][19] ) );
  DFFARX1 \FIFO_reg[13][18]  ( .D(n4133), .CLK(clk_in), .RSTB(n7130), .Q(
        \FIFO[13][18] ) );
  DFFARX1 \FIFO_reg[13][17]  ( .D(n4132), .CLK(clk_in), .RSTB(n7130), .Q(
        \FIFO[13][17] ) );
  DFFARX1 \FIFO_reg[13][16]  ( .D(n4131), .CLK(clk_in), .RSTB(n7130), .Q(
        \FIFO[13][16] ) );
  DFFARX1 \FIFO_reg[13][15]  ( .D(n4130), .CLK(clk_in), .RSTB(n7130), .Q(
        \FIFO[13][15] ) );
  DFFARX1 \FIFO_reg[13][14]  ( .D(n4129), .CLK(clk_in), .RSTB(n7130), .Q(
        \FIFO[13][14] ) );
  DFFARX1 \FIFO_reg[13][13]  ( .D(n4128), .CLK(clk_in), .RSTB(n7130), .Q(
        \FIFO[13][13] ) );
  DFFARX1 \FIFO_reg[13][12]  ( .D(n4127), .CLK(clk_in), .RSTB(n7130), .Q(
        \FIFO[13][12] ) );
  DFFARX1 \FIFO_reg[13][11]  ( .D(n4126), .CLK(clk_in), .RSTB(n7130), .Q(
        \FIFO[13][11] ) );
  DFFARX1 \FIFO_reg[13][10]  ( .D(n4125), .CLK(clk_in), .RSTB(n7130), .Q(
        \FIFO[13][10] ) );
  DFFARX1 \FIFO_reg[13][9]  ( .D(n4124), .CLK(clk_in), .RSTB(n7131), .Q(
        \FIFO[13][9] ) );
  DFFARX1 \FIFO_reg[13][8]  ( .D(n4123), .CLK(clk_in), .RSTB(n7131), .Q(
        \FIFO[13][8] ) );
  DFFARX1 \FIFO_reg[13][7]  ( .D(n4122), .CLK(clk_in), .RSTB(n7131), .Q(
        \FIFO[13][7] ) );
  DFFARX1 \FIFO_reg[13][6]  ( .D(n4121), .CLK(clk_in), .RSTB(n7131), .Q(
        \FIFO[13][6] ) );
  DFFARX1 \FIFO_reg[13][5]  ( .D(n4120), .CLK(clk_in), .RSTB(n7131), .Q(
        \FIFO[13][5] ) );
  DFFARX1 \FIFO_reg[13][4]  ( .D(n4119), .CLK(clk_in), .RSTB(n7131), .Q(
        \FIFO[13][4] ) );
  DFFARX1 \FIFO_reg[13][3]  ( .D(n4118), .CLK(clk_in), .RSTB(n7131), .Q(
        \FIFO[13][3] ) );
  DFFARX1 \FIFO_reg[13][2]  ( .D(n4117), .CLK(clk_in), .RSTB(n7131), .Q(
        \FIFO[13][2] ) );
  DFFARX1 \FIFO_reg[13][1]  ( .D(n4116), .CLK(clk_in), .RSTB(n7131), .Q(
        \FIFO[13][1] ) );
  DFFARX1 \FIFO_reg[13][0]  ( .D(n4115), .CLK(clk_in), .RSTB(n7131), .Q(
        \FIFO[13][0] ) );
  DFFARX1 \FIFO_reg[14][31]  ( .D(n4114), .CLK(clk_in), .RSTB(n7131), .Q(
        \FIFO[14][31] ) );
  DFFARX1 \FIFO_reg[14][30]  ( .D(n4113), .CLK(clk_in), .RSTB(n7131), .Q(
        \FIFO[14][30] ) );
  DFFARX1 \FIFO_reg[14][29]  ( .D(n4112), .CLK(clk_in), .RSTB(n7131), .Q(
        \FIFO[14][29] ) );
  DFFARX1 \FIFO_reg[14][28]  ( .D(n4111), .CLK(clk_in), .RSTB(n7131), .Q(
        \FIFO[14][28] ) );
  DFFARX1 \FIFO_reg[14][27]  ( .D(n4110), .CLK(clk_in), .RSTB(n7131), .Q(
        \FIFO[14][27] ) );
  DFFARX1 \FIFO_reg[14][26]  ( .D(n4109), .CLK(clk_in), .RSTB(n7131), .Q(
        \FIFO[14][26] ) );
  DFFARX1 \FIFO_reg[14][25]  ( .D(n4108), .CLK(clk_in), .RSTB(n7131), .Q(
        \FIFO[14][25] ) );
  DFFARX1 \FIFO_reg[14][24]  ( .D(n4107), .CLK(clk_in), .RSTB(n7131), .Q(
        \FIFO[14][24] ) );
  DFFARX1 \FIFO_reg[14][23]  ( .D(n4106), .CLK(clk_in), .RSTB(n7132), .Q(
        \FIFO[14][23] ) );
  DFFARX1 \FIFO_reg[14][22]  ( .D(n4105), .CLK(clk_in), .RSTB(n7132), .Q(
        \FIFO[14][22] ) );
  DFFARX1 \FIFO_reg[14][21]  ( .D(n4104), .CLK(clk_in), .RSTB(n7132), .Q(
        \FIFO[14][21] ) );
  DFFARX1 \FIFO_reg[14][20]  ( .D(n4103), .CLK(clk_in), .RSTB(n7132), .Q(
        \FIFO[14][20] ) );
  DFFARX1 \FIFO_reg[14][19]  ( .D(n4102), .CLK(clk_in), .RSTB(n7132), .Q(
        \FIFO[14][19] ) );
  DFFARX1 \FIFO_reg[14][18]  ( .D(n4101), .CLK(clk_in), .RSTB(n7132), .Q(
        \FIFO[14][18] ) );
  DFFARX1 \FIFO_reg[14][17]  ( .D(n4100), .CLK(clk_in), .RSTB(n7132), .Q(
        \FIFO[14][17] ) );
  DFFARX1 \FIFO_reg[14][16]  ( .D(n4099), .CLK(clk_in), .RSTB(n7132), .Q(
        \FIFO[14][16] ) );
  DFFARX1 \FIFO_reg[14][15]  ( .D(n4098), .CLK(clk_in), .RSTB(n7132), .Q(
        \FIFO[14][15] ) );
  DFFARX1 \FIFO_reg[14][14]  ( .D(n4097), .CLK(clk_in), .RSTB(n7132), .Q(
        \FIFO[14][14] ) );
  DFFARX1 \FIFO_reg[14][13]  ( .D(n4096), .CLK(clk_in), .RSTB(n7132), .Q(
        \FIFO[14][13] ) );
  DFFARX1 \FIFO_reg[14][12]  ( .D(n4095), .CLK(clk_in), .RSTB(n7132), .Q(
        \FIFO[14][12] ) );
  DFFARX1 \FIFO_reg[14][11]  ( .D(n4094), .CLK(clk_in), .RSTB(n7132), .Q(
        \FIFO[14][11] ) );
  DFFARX1 \FIFO_reg[14][10]  ( .D(n4093), .CLK(clk_in), .RSTB(n7132), .Q(
        \FIFO[14][10] ) );
  DFFARX1 \FIFO_reg[14][9]  ( .D(n4092), .CLK(clk_in), .RSTB(n7132), .Q(
        \FIFO[14][9] ) );
  DFFARX1 \FIFO_reg[14][8]  ( .D(n4091), .CLK(clk_in), .RSTB(n7132), .Q(
        \FIFO[14][8] ) );
  DFFARX1 \FIFO_reg[14][7]  ( .D(n4090), .CLK(clk_in), .RSTB(n7132), .Q(
        \FIFO[14][7] ) );
  DFFARX1 \FIFO_reg[14][6]  ( .D(n4089), .CLK(clk_in), .RSTB(n7132), .Q(
        \FIFO[14][6] ) );
  DFFARX1 \FIFO_reg[14][5]  ( .D(n4088), .CLK(clk_in), .RSTB(n7133), .Q(
        \FIFO[14][5] ) );
  DFFARX1 \FIFO_reg[14][4]  ( .D(n4087), .CLK(clk_in), .RSTB(n7133), .Q(
        \FIFO[14][4] ) );
  DFFARX1 \FIFO_reg[14][3]  ( .D(n4086), .CLK(clk_in), .RSTB(n7133), .Q(
        \FIFO[14][3] ) );
  DFFARX1 \FIFO_reg[14][2]  ( .D(n4085), .CLK(clk_in), .RSTB(n7133), .Q(
        \FIFO[14][2] ) );
  DFFARX1 \FIFO_reg[14][1]  ( .D(n4084), .CLK(clk_in), .RSTB(n7133), .Q(
        \FIFO[14][1] ) );
  DFFARX1 \FIFO_reg[14][0]  ( .D(n4083), .CLK(clk_in), .RSTB(n7133), .Q(
        \FIFO[14][0] ) );
  DFFARX1 \FIFO_reg[15][31]  ( .D(n4082), .CLK(clk_in), .RSTB(n7133), .Q(
        \FIFO[15][31] ) );
  DFFARX1 \FIFO_reg[15][30]  ( .D(n4081), .CLK(clk_in), .RSTB(n7133), .Q(
        \FIFO[15][30] ) );
  DFFARX1 \FIFO_reg[15][29]  ( .D(n4080), .CLK(clk_in), .RSTB(n7133), .Q(
        \FIFO[15][29] ) );
  DFFARX1 \FIFO_reg[15][28]  ( .D(n4079), .CLK(clk_in), .RSTB(n7133), .Q(
        \FIFO[15][28] ) );
  DFFARX1 \FIFO_reg[15][27]  ( .D(n4078), .CLK(clk_in), .RSTB(n7133), .Q(
        \FIFO[15][27] ) );
  DFFARX1 \FIFO_reg[15][26]  ( .D(n4077), .CLK(clk_in), .RSTB(n7133), .Q(
        \FIFO[15][26] ) );
  DFFARX1 \FIFO_reg[15][25]  ( .D(n4076), .CLK(clk_in), .RSTB(n7133), .Q(
        \FIFO[15][25] ) );
  DFFARX1 \FIFO_reg[15][24]  ( .D(n4075), .CLK(clk_in), .RSTB(n7133), .Q(
        \FIFO[15][24] ) );
  DFFARX1 \FIFO_reg[15][23]  ( .D(n4074), .CLK(clk_in), .RSTB(n7133), .Q(
        \FIFO[15][23] ) );
  DFFARX1 \FIFO_reg[15][22]  ( .D(n4073), .CLK(clk_in), .RSTB(n7133), .Q(
        \FIFO[15][22] ) );
  DFFARX1 \FIFO_reg[15][21]  ( .D(n4072), .CLK(clk_in), .RSTB(n7133), .Q(
        \FIFO[15][21] ) );
  DFFARX1 \FIFO_reg[15][20]  ( .D(n4071), .CLK(clk_in), .RSTB(n7133), .Q(
        \FIFO[15][20] ) );
  DFFARX1 \FIFO_reg[15][19]  ( .D(n4070), .CLK(clk_in), .RSTB(n7134), .Q(
        \FIFO[15][19] ) );
  DFFARX1 \FIFO_reg[15][18]  ( .D(n4069), .CLK(clk_in), .RSTB(n7134), .Q(
        \FIFO[15][18] ) );
  DFFARX1 \FIFO_reg[15][17]  ( .D(n4068), .CLK(clk_in), .RSTB(n7134), .Q(
        \FIFO[15][17] ) );
  DFFARX1 \FIFO_reg[15][16]  ( .D(n4067), .CLK(clk_in), .RSTB(n7134), .Q(
        \FIFO[15][16] ) );
  DFFARX1 \FIFO_reg[15][15]  ( .D(n4066), .CLK(clk_in), .RSTB(n7134), .Q(
        \FIFO[15][15] ) );
  DFFARX1 \FIFO_reg[15][14]  ( .D(n4065), .CLK(clk_in), .RSTB(n7134), .Q(
        \FIFO[15][14] ) );
  DFFARX1 \FIFO_reg[15][13]  ( .D(n4064), .CLK(clk_in), .RSTB(n7134), .Q(
        \FIFO[15][13] ) );
  DFFARX1 \FIFO_reg[15][12]  ( .D(n4063), .CLK(clk_in), .RSTB(n7134), .Q(
        \FIFO[15][12] ) );
  DFFARX1 \FIFO_reg[15][11]  ( .D(n4062), .CLK(clk_in), .RSTB(n7134), .Q(
        \FIFO[15][11] ) );
  DFFARX1 \FIFO_reg[15][10]  ( .D(n4061), .CLK(clk_in), .RSTB(n7134), .Q(
        \FIFO[15][10] ) );
  DFFARX1 \FIFO_reg[15][9]  ( .D(n4060), .CLK(clk_in), .RSTB(n7134), .Q(
        \FIFO[15][9] ) );
  DFFARX1 \FIFO_reg[15][8]  ( .D(n4059), .CLK(clk_in), .RSTB(n7134), .Q(
        \FIFO[15][8] ) );
  DFFARX1 \FIFO_reg[15][7]  ( .D(n4058), .CLK(clk_in), .RSTB(n7134), .Q(
        \FIFO[15][7] ) );
  DFFARX1 \FIFO_reg[15][6]  ( .D(n4057), .CLK(clk_in), .RSTB(n7134), .Q(
        \FIFO[15][6] ) );
  DFFARX1 \FIFO_reg[15][5]  ( .D(n4056), .CLK(clk_in), .RSTB(n7134), .Q(
        \FIFO[15][5] ) );
  DFFARX1 \FIFO_reg[15][4]  ( .D(n4055), .CLK(clk_in), .RSTB(n7134), .Q(
        \FIFO[15][4] ) );
  DFFARX1 \FIFO_reg[15][3]  ( .D(n4054), .CLK(clk_in), .RSTB(n7134), .Q(
        \FIFO[15][3] ) );
  DFFARX1 \FIFO_reg[15][2]  ( .D(n4053), .CLK(clk_in), .RSTB(n7134), .Q(
        \FIFO[15][2] ) );
  DFFARX1 \FIFO_reg[15][1]  ( .D(n4052), .CLK(clk_in), .RSTB(n7135), .Q(
        \FIFO[15][1] ) );
  DFFARX1 \FIFO_reg[15][0]  ( .D(n4051), .CLK(clk_in), .RSTB(n7135), .Q(
        \FIFO[15][0] ) );
  DFFARX1 \FIFO_reg[16][31]  ( .D(n4050), .CLK(clk_in), .RSTB(n7135), .Q(
        \FIFO[16][31] ) );
  DFFARX1 \FIFO_reg[16][30]  ( .D(n4049), .CLK(clk_in), .RSTB(n7135), .Q(
        \FIFO[16][30] ) );
  DFFARX1 \FIFO_reg[16][29]  ( .D(n4048), .CLK(clk_in), .RSTB(n7135), .Q(
        \FIFO[16][29] ) );
  DFFARX1 \FIFO_reg[16][28]  ( .D(n4047), .CLK(clk_in), .RSTB(n7135), .Q(
        \FIFO[16][28] ) );
  DFFARX1 \FIFO_reg[16][27]  ( .D(n4046), .CLK(clk_in), .RSTB(n7135), .Q(
        \FIFO[16][27] ) );
  DFFARX1 \FIFO_reg[16][26]  ( .D(n4045), .CLK(clk_in), .RSTB(n7135), .Q(
        \FIFO[16][26] ) );
  DFFARX1 \FIFO_reg[16][25]  ( .D(n4044), .CLK(clk_in), .RSTB(n7135), .Q(
        \FIFO[16][25] ) );
  DFFARX1 \FIFO_reg[16][24]  ( .D(n4043), .CLK(clk_in), .RSTB(n7135), .Q(
        \FIFO[16][24] ) );
  DFFARX1 \FIFO_reg[16][23]  ( .D(n4042), .CLK(clk_in), .RSTB(n7135), .Q(
        \FIFO[16][23] ) );
  DFFARX1 \FIFO_reg[16][22]  ( .D(n4041), .CLK(clk_in), .RSTB(n7135), .Q(
        \FIFO[16][22] ) );
  DFFARX1 \FIFO_reg[16][21]  ( .D(n4040), .CLK(clk_in), .RSTB(n7135), .Q(
        \FIFO[16][21] ) );
  DFFARX1 \FIFO_reg[16][20]  ( .D(n4039), .CLK(clk_in), .RSTB(n7135), .Q(
        \FIFO[16][20] ) );
  DFFARX1 \FIFO_reg[16][19]  ( .D(n4038), .CLK(clk_in), .RSTB(n7135), .Q(
        \FIFO[16][19] ) );
  DFFARX1 \FIFO_reg[16][18]  ( .D(n4037), .CLK(clk_in), .RSTB(n7135), .Q(
        \FIFO[16][18] ) );
  DFFARX1 \FIFO_reg[16][17]  ( .D(n4036), .CLK(clk_in), .RSTB(n7135), .Q(
        \FIFO[16][17] ) );
  DFFARX1 \FIFO_reg[16][16]  ( .D(n4035), .CLK(clk_in), .RSTB(n7135), .Q(
        \FIFO[16][16] ) );
  DFFARX1 \FIFO_reg[16][15]  ( .D(n4034), .CLK(clk_in), .RSTB(n7136), .Q(
        \FIFO[16][15] ) );
  DFFARX1 \FIFO_reg[16][14]  ( .D(n4033), .CLK(clk_in), .RSTB(n7136), .Q(
        \FIFO[16][14] ) );
  DFFARX1 \FIFO_reg[16][13]  ( .D(n4032), .CLK(clk_in), .RSTB(n7136), .Q(
        \FIFO[16][13] ) );
  DFFARX1 \FIFO_reg[16][12]  ( .D(n4031), .CLK(clk_in), .RSTB(n7136), .Q(
        \FIFO[16][12] ) );
  DFFARX1 \FIFO_reg[16][11]  ( .D(n4030), .CLK(clk_in), .RSTB(n7136), .Q(
        \FIFO[16][11] ) );
  DFFARX1 \FIFO_reg[16][10]  ( .D(n4029), .CLK(clk_in), .RSTB(n7136), .Q(
        \FIFO[16][10] ) );
  DFFARX1 \FIFO_reg[16][9]  ( .D(n4028), .CLK(clk_in), .RSTB(n7136), .Q(
        \FIFO[16][9] ) );
  DFFARX1 \FIFO_reg[16][8]  ( .D(n4027), .CLK(clk_in), .RSTB(n7136), .Q(
        \FIFO[16][8] ) );
  DFFARX1 \FIFO_reg[16][7]  ( .D(n4026), .CLK(clk_in), .RSTB(n7136), .Q(
        \FIFO[16][7] ) );
  DFFARX1 \FIFO_reg[16][6]  ( .D(n4025), .CLK(clk_in), .RSTB(n7136), .Q(
        \FIFO[16][6] ) );
  DFFARX1 \FIFO_reg[16][5]  ( .D(n4024), .CLK(clk_in), .RSTB(n7136), .Q(
        \FIFO[16][5] ) );
  DFFARX1 \FIFO_reg[16][4]  ( .D(n4023), .CLK(clk_in), .RSTB(n7136), .Q(
        \FIFO[16][4] ) );
  DFFARX1 \FIFO_reg[16][3]  ( .D(n4022), .CLK(clk_in), .RSTB(n7136), .Q(
        \FIFO[16][3] ) );
  DFFARX1 \FIFO_reg[16][2]  ( .D(n4021), .CLK(clk_in), .RSTB(n7136), .Q(
        \FIFO[16][2] ) );
  DFFARX1 \FIFO_reg[16][1]  ( .D(n4020), .CLK(clk_in), .RSTB(n7136), .Q(
        \FIFO[16][1] ) );
  DFFARX1 \FIFO_reg[16][0]  ( .D(n4019), .CLK(clk_in), .RSTB(n7136), .Q(
        \FIFO[16][0] ) );
  DFFARX1 \FIFO_reg[17][31]  ( .D(n4018), .CLK(clk_in), .RSTB(n7136), .Q(
        \FIFO[17][31] ) );
  DFFARX1 \FIFO_reg[17][30]  ( .D(n4017), .CLK(clk_in), .RSTB(n7136), .Q(
        \FIFO[17][30] ) );
  DFFARX1 \FIFO_reg[17][29]  ( .D(n4016), .CLK(clk_in), .RSTB(n7137), .Q(
        \FIFO[17][29] ) );
  DFFARX1 \FIFO_reg[17][28]  ( .D(n4015), .CLK(clk_in), .RSTB(n7137), .Q(
        \FIFO[17][28] ) );
  DFFARX1 \FIFO_reg[17][27]  ( .D(n4014), .CLK(clk_in), .RSTB(n7137), .Q(
        \FIFO[17][27] ) );
  DFFARX1 \FIFO_reg[17][26]  ( .D(n4013), .CLK(clk_in), .RSTB(n7137), .Q(
        \FIFO[17][26] ) );
  DFFARX1 \FIFO_reg[17][25]  ( .D(n4012), .CLK(clk_in), .RSTB(n7137), .Q(
        \FIFO[17][25] ) );
  DFFARX1 \FIFO_reg[17][24]  ( .D(n4011), .CLK(clk_in), .RSTB(n7137), .Q(
        \FIFO[17][24] ) );
  DFFARX1 \FIFO_reg[17][23]  ( .D(n4010), .CLK(clk_in), .RSTB(n7137), .Q(
        \FIFO[17][23] ) );
  DFFARX1 \FIFO_reg[17][22]  ( .D(n4009), .CLK(clk_in), .RSTB(n7137), .Q(
        \FIFO[17][22] ) );
  DFFARX1 \FIFO_reg[17][21]  ( .D(n4008), .CLK(clk_in), .RSTB(n7137), .Q(
        \FIFO[17][21] ) );
  DFFARX1 \FIFO_reg[17][20]  ( .D(n4007), .CLK(clk_in), .RSTB(n7137), .Q(
        \FIFO[17][20] ) );
  DFFARX1 \FIFO_reg[17][19]  ( .D(n4006), .CLK(clk_in), .RSTB(n7137), .Q(
        \FIFO[17][19] ) );
  DFFARX1 \FIFO_reg[17][18]  ( .D(n4005), .CLK(clk_in), .RSTB(n7137), .Q(
        \FIFO[17][18] ) );
  DFFARX1 \FIFO_reg[17][17]  ( .D(n4004), .CLK(clk_in), .RSTB(n7137), .Q(
        \FIFO[17][17] ) );
  DFFARX1 \FIFO_reg[17][16]  ( .D(n4003), .CLK(clk_in), .RSTB(n7137), .Q(
        \FIFO[17][16] ) );
  DFFARX1 \FIFO_reg[17][15]  ( .D(n4002), .CLK(clk_in), .RSTB(n7137), .Q(
        \FIFO[17][15] ) );
  DFFARX1 \FIFO_reg[17][14]  ( .D(n4001), .CLK(clk_in), .RSTB(n7137), .Q(
        \FIFO[17][14] ) );
  DFFARX1 \FIFO_reg[17][13]  ( .D(n4000), .CLK(clk_in), .RSTB(n7137), .Q(
        \FIFO[17][13] ) );
  DFFARX1 \FIFO_reg[17][12]  ( .D(n3999), .CLK(clk_in), .RSTB(n7137), .Q(
        \FIFO[17][12] ) );
  DFFARX1 \FIFO_reg[17][11]  ( .D(n3998), .CLK(clk_in), .RSTB(n7138), .Q(
        \FIFO[17][11] ) );
  DFFARX1 \FIFO_reg[17][10]  ( .D(n3997), .CLK(clk_in), .RSTB(n7138), .Q(
        \FIFO[17][10] ) );
  DFFARX1 \FIFO_reg[17][9]  ( .D(n3996), .CLK(clk_in), .RSTB(n7138), .Q(
        \FIFO[17][9] ) );
  DFFARX1 \FIFO_reg[17][8]  ( .D(n3995), .CLK(clk_in), .RSTB(n7138), .Q(
        \FIFO[17][8] ) );
  DFFARX1 \FIFO_reg[17][7]  ( .D(n3994), .CLK(clk_in), .RSTB(n7138), .Q(
        \FIFO[17][7] ) );
  DFFARX1 \FIFO_reg[17][6]  ( .D(n3993), .CLK(clk_in), .RSTB(n7138), .Q(
        \FIFO[17][6] ) );
  DFFARX1 \FIFO_reg[17][5]  ( .D(n3992), .CLK(clk_in), .RSTB(n7138), .Q(
        \FIFO[17][5] ) );
  DFFARX1 \FIFO_reg[17][4]  ( .D(n3991), .CLK(clk_in), .RSTB(n7138), .Q(
        \FIFO[17][4] ) );
  DFFARX1 \FIFO_reg[17][3]  ( .D(n3990), .CLK(clk_in), .RSTB(n7138), .Q(
        \FIFO[17][3] ) );
  DFFARX1 \FIFO_reg[17][2]  ( .D(n3989), .CLK(clk_in), .RSTB(n7138), .Q(
        \FIFO[17][2] ) );
  DFFARX1 \FIFO_reg[17][1]  ( .D(n3988), .CLK(clk_in), .RSTB(n7138), .Q(
        \FIFO[17][1] ) );
  DFFARX1 \FIFO_reg[17][0]  ( .D(n3987), .CLK(clk_in), .RSTB(n7138), .Q(
        \FIFO[17][0] ) );
  DFFARX1 \FIFO_reg[18][31]  ( .D(n3986), .CLK(clk_in), .RSTB(n7138), .Q(
        \FIFO[18][31] ) );
  DFFARX1 \FIFO_reg[18][30]  ( .D(n3985), .CLK(clk_in), .RSTB(n7138), .Q(
        \FIFO[18][30] ) );
  DFFARX1 \FIFO_reg[18][29]  ( .D(n3984), .CLK(clk_in), .RSTB(n7138), .Q(
        \FIFO[18][29] ) );
  DFFARX1 \FIFO_reg[18][28]  ( .D(n3983), .CLK(clk_in), .RSTB(n7138), .Q(
        \FIFO[18][28] ) );
  DFFARX1 \FIFO_reg[18][27]  ( .D(n3982), .CLK(clk_in), .RSTB(n7138), .Q(
        \FIFO[18][27] ) );
  DFFARX1 \FIFO_reg[18][26]  ( .D(n3981), .CLK(clk_in), .RSTB(n7138), .Q(
        \FIFO[18][26] ) );
  DFFARX1 \FIFO_reg[18][25]  ( .D(n3980), .CLK(clk_in), .RSTB(n7139), .Q(
        \FIFO[18][25] ) );
  DFFARX1 \FIFO_reg[18][24]  ( .D(n3979), .CLK(clk_in), .RSTB(n7139), .Q(
        \FIFO[18][24] ) );
  DFFARX1 \FIFO_reg[18][23]  ( .D(n3978), .CLK(clk_in), .RSTB(n7139), .Q(
        \FIFO[18][23] ) );
  DFFARX1 \FIFO_reg[18][22]  ( .D(n3977), .CLK(clk_in), .RSTB(n7139), .Q(
        \FIFO[18][22] ) );
  DFFARX1 \FIFO_reg[18][21]  ( .D(n3976), .CLK(clk_in), .RSTB(n7139), .Q(
        \FIFO[18][21] ) );
  DFFARX1 \FIFO_reg[18][20]  ( .D(n3975), .CLK(clk_in), .RSTB(n7139), .Q(
        \FIFO[18][20] ) );
  DFFARX1 \FIFO_reg[18][19]  ( .D(n3974), .CLK(clk_in), .RSTB(n7139), .Q(
        \FIFO[18][19] ) );
  DFFARX1 \FIFO_reg[18][18]  ( .D(n3973), .CLK(clk_in), .RSTB(n7139), .Q(
        \FIFO[18][18] ) );
  DFFARX1 \FIFO_reg[18][17]  ( .D(n3972), .CLK(clk_in), .RSTB(n7139), .Q(
        \FIFO[18][17] ) );
  DFFARX1 \FIFO_reg[18][16]  ( .D(n3971), .CLK(clk_in), .RSTB(n7139), .Q(
        \FIFO[18][16] ) );
  DFFARX1 \FIFO_reg[18][15]  ( .D(n3970), .CLK(clk_in), .RSTB(n7139), .Q(
        \FIFO[18][15] ) );
  DFFARX1 \FIFO_reg[18][14]  ( .D(n3969), .CLK(clk_in), .RSTB(n7139), .Q(
        \FIFO[18][14] ) );
  DFFARX1 \FIFO_reg[18][13]  ( .D(n3968), .CLK(clk_in), .RSTB(n7139), .Q(
        \FIFO[18][13] ) );
  DFFARX1 \FIFO_reg[18][12]  ( .D(n3967), .CLK(clk_in), .RSTB(n7139), .Q(
        \FIFO[18][12] ) );
  DFFARX1 \FIFO_reg[18][11]  ( .D(n3966), .CLK(clk_in), .RSTB(n7139), .Q(
        \FIFO[18][11] ) );
  DFFARX1 \FIFO_reg[18][10]  ( .D(n3965), .CLK(clk_in), .RSTB(n7139), .Q(
        \FIFO[18][10] ) );
  DFFARX1 \FIFO_reg[18][9]  ( .D(n3964), .CLK(clk_in), .RSTB(n7139), .Q(
        \FIFO[18][9] ) );
  DFFARX1 \FIFO_reg[18][8]  ( .D(n3963), .CLK(clk_in), .RSTB(n7139), .Q(
        \FIFO[18][8] ) );
  DFFARX1 \FIFO_reg[18][7]  ( .D(n3962), .CLK(clk_in), .RSTB(n7140), .Q(
        \FIFO[18][7] ) );
  DFFARX1 \FIFO_reg[18][6]  ( .D(n3961), .CLK(clk_in), .RSTB(n7140), .Q(
        \FIFO[18][6] ) );
  DFFARX1 \FIFO_reg[18][5]  ( .D(n3960), .CLK(clk_in), .RSTB(n7140), .Q(
        \FIFO[18][5] ) );
  DFFARX1 \FIFO_reg[18][4]  ( .D(n3959), .CLK(clk_in), .RSTB(n7140), .Q(
        \FIFO[18][4] ) );
  DFFARX1 \FIFO_reg[18][3]  ( .D(n3958), .CLK(clk_in), .RSTB(n7140), .Q(
        \FIFO[18][3] ) );
  DFFARX1 \FIFO_reg[18][2]  ( .D(n3957), .CLK(clk_in), .RSTB(n7140), .Q(
        \FIFO[18][2] ) );
  DFFARX1 \FIFO_reg[18][1]  ( .D(n3956), .CLK(clk_in), .RSTB(n7140), .Q(
        \FIFO[18][1] ) );
  DFFARX1 \FIFO_reg[18][0]  ( .D(n3955), .CLK(clk_in), .RSTB(n7140), .Q(
        \FIFO[18][0] ) );
  DFFARX1 \FIFO_reg[19][31]  ( .D(n3954), .CLK(clk_in), .RSTB(n7140), .Q(
        \FIFO[19][31] ) );
  DFFARX1 \FIFO_reg[19][30]  ( .D(n3953), .CLK(clk_in), .RSTB(n7140), .Q(
        \FIFO[19][30] ) );
  DFFARX1 \FIFO_reg[19][29]  ( .D(n3952), .CLK(clk_in), .RSTB(n7140), .Q(
        \FIFO[19][29] ) );
  DFFARX1 \FIFO_reg[19][28]  ( .D(n3951), .CLK(clk_in), .RSTB(n7140), .Q(
        \FIFO[19][28] ) );
  DFFARX1 \FIFO_reg[19][27]  ( .D(n3950), .CLK(clk_in), .RSTB(n7140), .Q(
        \FIFO[19][27] ) );
  DFFARX1 \FIFO_reg[19][26]  ( .D(n3949), .CLK(clk_in), .RSTB(n7140), .Q(
        \FIFO[19][26] ) );
  DFFARX1 \FIFO_reg[19][25]  ( .D(n3948), .CLK(clk_in), .RSTB(n7140), .Q(
        \FIFO[19][25] ) );
  DFFARX1 \FIFO_reg[19][24]  ( .D(n3947), .CLK(clk_in), .RSTB(n7140), .Q(
        \FIFO[19][24] ) );
  DFFARX1 \FIFO_reg[19][23]  ( .D(n3946), .CLK(clk_in), .RSTB(n7140), .Q(
        \FIFO[19][23] ) );
  DFFARX1 \FIFO_reg[19][22]  ( .D(n3945), .CLK(clk_in), .RSTB(n7140), .Q(
        \FIFO[19][22] ) );
  DFFARX1 \FIFO_reg[19][21]  ( .D(n3944), .CLK(clk_in), .RSTB(n7141), .Q(
        \FIFO[19][21] ) );
  DFFARX1 \FIFO_reg[19][20]  ( .D(n3943), .CLK(clk_in), .RSTB(n7141), .Q(
        \FIFO[19][20] ) );
  DFFARX1 \FIFO_reg[19][19]  ( .D(n3942), .CLK(clk_in), .RSTB(n7141), .Q(
        \FIFO[19][19] ) );
  DFFARX1 \FIFO_reg[19][18]  ( .D(n3941), .CLK(clk_in), .RSTB(n7141), .Q(
        \FIFO[19][18] ) );
  DFFARX1 \FIFO_reg[19][17]  ( .D(n3940), .CLK(clk_in), .RSTB(n7141), .Q(
        \FIFO[19][17] ) );
  DFFARX1 \FIFO_reg[19][16]  ( .D(n3939), .CLK(clk_in), .RSTB(n7141), .Q(
        \FIFO[19][16] ) );
  DFFARX1 \FIFO_reg[19][15]  ( .D(n3938), .CLK(clk_in), .RSTB(n7141), .Q(
        \FIFO[19][15] ) );
  DFFARX1 \FIFO_reg[19][14]  ( .D(n3937), .CLK(clk_in), .RSTB(n7141), .Q(
        \FIFO[19][14] ) );
  DFFARX1 \FIFO_reg[19][13]  ( .D(n3936), .CLK(clk_in), .RSTB(n7141), .Q(
        \FIFO[19][13] ) );
  DFFARX1 \FIFO_reg[19][12]  ( .D(n3935), .CLK(clk_in), .RSTB(n7141), .Q(
        \FIFO[19][12] ) );
  DFFARX1 \FIFO_reg[19][11]  ( .D(n3934), .CLK(clk_in), .RSTB(n7141), .Q(
        \FIFO[19][11] ) );
  DFFARX1 \FIFO_reg[19][10]  ( .D(n3933), .CLK(clk_in), .RSTB(n7141), .Q(
        \FIFO[19][10] ) );
  DFFARX1 \FIFO_reg[19][9]  ( .D(n3932), .CLK(clk_in), .RSTB(n7141), .Q(
        \FIFO[19][9] ) );
  DFFARX1 \FIFO_reg[19][8]  ( .D(n3931), .CLK(clk_in), .RSTB(n7141), .Q(
        \FIFO[19][8] ) );
  DFFARX1 \FIFO_reg[19][7]  ( .D(n3930), .CLK(clk_in), .RSTB(n7141), .Q(
        \FIFO[19][7] ) );
  DFFARX1 \FIFO_reg[19][6]  ( .D(n3929), .CLK(clk_in), .RSTB(n7141), .Q(
        \FIFO[19][6] ) );
  DFFARX1 \FIFO_reg[19][5]  ( .D(n3928), .CLK(clk_in), .RSTB(n7141), .Q(
        \FIFO[19][5] ) );
  DFFARX1 \FIFO_reg[19][4]  ( .D(n3927), .CLK(clk_in), .RSTB(n7141), .Q(
        \FIFO[19][4] ) );
  DFFARX1 \FIFO_reg[19][3]  ( .D(n3926), .CLK(clk_in), .RSTB(n7142), .Q(
        \FIFO[19][3] ) );
  DFFARX1 \FIFO_reg[19][2]  ( .D(n3925), .CLK(clk_in), .RSTB(n7142), .Q(
        \FIFO[19][2] ) );
  DFFARX1 \FIFO_reg[19][1]  ( .D(n3924), .CLK(clk_in), .RSTB(n7142), .Q(
        \FIFO[19][1] ) );
  DFFARX1 \FIFO_reg[19][0]  ( .D(n3923), .CLK(clk_in), .RSTB(n7142), .Q(
        \FIFO[19][0] ) );
  DFFARX1 \FIFO_reg[20][31]  ( .D(n3922), .CLK(clk_in), .RSTB(n7142), .Q(
        \FIFO[20][31] ) );
  DFFARX1 \FIFO_reg[20][30]  ( .D(n3921), .CLK(clk_in), .RSTB(n7142), .Q(
        \FIFO[20][30] ) );
  DFFARX1 \FIFO_reg[20][29]  ( .D(n3920), .CLK(clk_in), .RSTB(n7142), .Q(
        \FIFO[20][29] ) );
  DFFARX1 \FIFO_reg[20][28]  ( .D(n3919), .CLK(clk_in), .RSTB(n7142), .Q(
        \FIFO[20][28] ) );
  DFFARX1 \FIFO_reg[20][27]  ( .D(n3918), .CLK(clk_in), .RSTB(n7142), .Q(
        \FIFO[20][27] ) );
  DFFARX1 \FIFO_reg[20][26]  ( .D(n3917), .CLK(clk_in), .RSTB(n7142), .Q(
        \FIFO[20][26] ) );
  DFFARX1 \FIFO_reg[20][25]  ( .D(n3916), .CLK(clk_in), .RSTB(n7142), .Q(
        \FIFO[20][25] ) );
  DFFARX1 \FIFO_reg[20][24]  ( .D(n3915), .CLK(clk_in), .RSTB(n7142), .Q(
        \FIFO[20][24] ) );
  DFFARX1 \FIFO_reg[20][23]  ( .D(n3914), .CLK(clk_in), .RSTB(n7142), .Q(
        \FIFO[20][23] ) );
  DFFARX1 \FIFO_reg[20][22]  ( .D(n3913), .CLK(clk_in), .RSTB(n7142), .Q(
        \FIFO[20][22] ) );
  DFFARX1 \FIFO_reg[20][21]  ( .D(n3912), .CLK(clk_in), .RSTB(n7142), .Q(
        \FIFO[20][21] ) );
  DFFARX1 \FIFO_reg[20][20]  ( .D(n3911), .CLK(clk_in), .RSTB(n7142), .Q(
        \FIFO[20][20] ) );
  DFFARX1 \FIFO_reg[20][19]  ( .D(n3910), .CLK(clk_in), .RSTB(n7142), .Q(
        \FIFO[20][19] ) );
  DFFARX1 \FIFO_reg[20][18]  ( .D(n3909), .CLK(clk_in), .RSTB(n7142), .Q(
        \FIFO[20][18] ) );
  DFFARX1 \FIFO_reg[20][17]  ( .D(n3908), .CLK(clk_in), .RSTB(n7143), .Q(
        \FIFO[20][17] ) );
  DFFARX1 \FIFO_reg[20][16]  ( .D(n3907), .CLK(clk_in), .RSTB(n7143), .Q(
        \FIFO[20][16] ) );
  DFFARX1 \FIFO_reg[20][15]  ( .D(n3906), .CLK(clk_in), .RSTB(n7143), .Q(
        \FIFO[20][15] ) );
  DFFARX1 \FIFO_reg[20][14]  ( .D(n3905), .CLK(clk_in), .RSTB(n7143), .Q(
        \FIFO[20][14] ) );
  DFFARX1 \FIFO_reg[20][13]  ( .D(n3904), .CLK(clk_in), .RSTB(n7143), .Q(
        \FIFO[20][13] ) );
  DFFARX1 \FIFO_reg[20][12]  ( .D(n3903), .CLK(clk_in), .RSTB(n7143), .Q(
        \FIFO[20][12] ) );
  DFFARX1 \FIFO_reg[20][11]  ( .D(n3902), .CLK(clk_in), .RSTB(n7143), .Q(
        \FIFO[20][11] ) );
  DFFARX1 \FIFO_reg[20][10]  ( .D(n3901), .CLK(clk_in), .RSTB(n7143), .Q(
        \FIFO[20][10] ) );
  DFFARX1 \FIFO_reg[20][9]  ( .D(n3900), .CLK(clk_in), .RSTB(n7143), .Q(
        \FIFO[20][9] ) );
  DFFARX1 \FIFO_reg[20][8]  ( .D(n3899), .CLK(clk_in), .RSTB(n7143), .Q(
        \FIFO[20][8] ) );
  DFFARX1 \FIFO_reg[20][7]  ( .D(n3898), .CLK(clk_in), .RSTB(n7143), .Q(
        \FIFO[20][7] ) );
  DFFARX1 \FIFO_reg[20][6]  ( .D(n3897), .CLK(clk_in), .RSTB(n7143), .Q(
        \FIFO[20][6] ) );
  DFFARX1 \FIFO_reg[20][5]  ( .D(n3896), .CLK(clk_in), .RSTB(n7143), .Q(
        \FIFO[20][5] ) );
  DFFARX1 \FIFO_reg[20][4]  ( .D(n3895), .CLK(clk_in), .RSTB(n7143), .Q(
        \FIFO[20][4] ) );
  DFFARX1 \FIFO_reg[20][3]  ( .D(n3894), .CLK(clk_in), .RSTB(n7143), .Q(
        \FIFO[20][3] ) );
  DFFARX1 \FIFO_reg[20][2]  ( .D(n3893), .CLK(clk_in), .RSTB(n7143), .Q(
        \FIFO[20][2] ) );
  DFFARX1 \FIFO_reg[20][1]  ( .D(n3892), .CLK(clk_in), .RSTB(n7143), .Q(
        \FIFO[20][1] ) );
  DFFARX1 \FIFO_reg[20][0]  ( .D(n3891), .CLK(clk_in), .RSTB(n7143), .Q(
        \FIFO[20][0] ) );
  DFFARX1 \FIFO_reg[21][31]  ( .D(n3890), .CLK(clk_in), .RSTB(n7144), .Q(
        \FIFO[21][31] ) );
  DFFARX1 \FIFO_reg[21][30]  ( .D(n3889), .CLK(clk_in), .RSTB(n7144), .Q(
        \FIFO[21][30] ) );
  DFFARX1 \FIFO_reg[21][29]  ( .D(n3888), .CLK(clk_in), .RSTB(n7144), .Q(
        \FIFO[21][29] ) );
  DFFARX1 \FIFO_reg[21][28]  ( .D(n3887), .CLK(clk_in), .RSTB(n7144), .Q(
        \FIFO[21][28] ) );
  DFFARX1 \FIFO_reg[21][27]  ( .D(n3886), .CLK(clk_in), .RSTB(n7144), .Q(
        \FIFO[21][27] ) );
  DFFARX1 \FIFO_reg[21][26]  ( .D(n3885), .CLK(clk_in), .RSTB(n7144), .Q(
        \FIFO[21][26] ) );
  DFFARX1 \FIFO_reg[21][25]  ( .D(n3884), .CLK(clk_in), .RSTB(n7144), .Q(
        \FIFO[21][25] ) );
  DFFARX1 \FIFO_reg[21][24]  ( .D(n3883), .CLK(clk_in), .RSTB(n7144), .Q(
        \FIFO[21][24] ) );
  DFFARX1 \FIFO_reg[21][23]  ( .D(n3882), .CLK(clk_in), .RSTB(n7144), .Q(
        \FIFO[21][23] ) );
  DFFARX1 \FIFO_reg[21][22]  ( .D(n3881), .CLK(clk_in), .RSTB(n7144), .Q(
        \FIFO[21][22] ) );
  DFFARX1 \FIFO_reg[21][21]  ( .D(n3880), .CLK(clk_in), .RSTB(n7144), .Q(
        \FIFO[21][21] ) );
  DFFARX1 \FIFO_reg[21][20]  ( .D(n3879), .CLK(clk_in), .RSTB(n7144), .Q(
        \FIFO[21][20] ) );
  DFFARX1 \FIFO_reg[21][19]  ( .D(n3878), .CLK(clk_in), .RSTB(n7144), .Q(
        \FIFO[21][19] ) );
  DFFARX1 \FIFO_reg[21][18]  ( .D(n3877), .CLK(clk_in), .RSTB(n7144), .Q(
        \FIFO[21][18] ) );
  DFFARX1 \FIFO_reg[21][17]  ( .D(n3876), .CLK(clk_in), .RSTB(n7144), .Q(
        \FIFO[21][17] ) );
  DFFARX1 \FIFO_reg[21][16]  ( .D(n3875), .CLK(clk_in), .RSTB(n7144), .Q(
        \FIFO[21][16] ) );
  DFFARX1 \FIFO_reg[21][15]  ( .D(n3874), .CLK(clk_in), .RSTB(n7144), .Q(
        \FIFO[21][15] ) );
  DFFARX1 \FIFO_reg[21][14]  ( .D(n3873), .CLK(clk_in), .RSTB(n7144), .Q(
        \FIFO[21][14] ) );
  DFFARX1 \FIFO_reg[21][13]  ( .D(n3872), .CLK(clk_in), .RSTB(n7145), .Q(
        \FIFO[21][13] ) );
  DFFARX1 \FIFO_reg[21][12]  ( .D(n3871), .CLK(clk_in), .RSTB(n7145), .Q(
        \FIFO[21][12] ) );
  DFFARX1 \FIFO_reg[21][11]  ( .D(n3870), .CLK(clk_in), .RSTB(n7145), .Q(
        \FIFO[21][11] ) );
  DFFARX1 \FIFO_reg[21][10]  ( .D(n3869), .CLK(clk_in), .RSTB(n7145), .Q(
        \FIFO[21][10] ) );
  DFFARX1 \FIFO_reg[21][9]  ( .D(n3868), .CLK(clk_in), .RSTB(n7145), .Q(
        \FIFO[21][9] ) );
  DFFARX1 \FIFO_reg[21][8]  ( .D(n3867), .CLK(clk_in), .RSTB(n7145), .Q(
        \FIFO[21][8] ) );
  DFFARX1 \FIFO_reg[21][7]  ( .D(n3866), .CLK(clk_in), .RSTB(n7145), .Q(
        \FIFO[21][7] ) );
  DFFARX1 \FIFO_reg[21][6]  ( .D(n3865), .CLK(clk_in), .RSTB(n7145), .Q(
        \FIFO[21][6] ) );
  DFFARX1 \FIFO_reg[21][5]  ( .D(n3864), .CLK(clk_in), .RSTB(n7145), .Q(
        \FIFO[21][5] ) );
  DFFARX1 \FIFO_reg[21][4]  ( .D(n3863), .CLK(clk_in), .RSTB(n7145), .Q(
        \FIFO[21][4] ) );
  DFFARX1 \FIFO_reg[21][3]  ( .D(n3862), .CLK(clk_in), .RSTB(n7145), .Q(
        \FIFO[21][3] ) );
  DFFARX1 \FIFO_reg[21][2]  ( .D(n3861), .CLK(clk_in), .RSTB(n7145), .Q(
        \FIFO[21][2] ) );
  DFFARX1 \FIFO_reg[21][1]  ( .D(n3860), .CLK(clk_in), .RSTB(n7145), .Q(
        \FIFO[21][1] ) );
  DFFARX1 \FIFO_reg[21][0]  ( .D(n3859), .CLK(clk_in), .RSTB(n7145), .Q(
        \FIFO[21][0] ) );
  DFFARX1 \FIFO_reg[22][31]  ( .D(n3858), .CLK(clk_in), .RSTB(n7145), .Q(
        \FIFO[22][31] ) );
  DFFARX1 \FIFO_reg[22][30]  ( .D(n3857), .CLK(clk_in), .RSTB(n7145), .Q(
        \FIFO[22][30] ) );
  DFFARX1 \FIFO_reg[22][29]  ( .D(n3856), .CLK(clk_in), .RSTB(n7145), .Q(
        \FIFO[22][29] ) );
  DFFARX1 \FIFO_reg[22][28]  ( .D(n3855), .CLK(clk_in), .RSTB(n7145), .Q(
        \FIFO[22][28] ) );
  DFFARX1 \FIFO_reg[22][27]  ( .D(n3854), .CLK(clk_in), .RSTB(n7146), .Q(
        \FIFO[22][27] ) );
  DFFARX1 \FIFO_reg[22][26]  ( .D(n3853), .CLK(clk_in), .RSTB(n7146), .Q(
        \FIFO[22][26] ) );
  DFFARX1 \FIFO_reg[22][25]  ( .D(n3852), .CLK(clk_in), .RSTB(n7146), .Q(
        \FIFO[22][25] ) );
  DFFARX1 \FIFO_reg[22][24]  ( .D(n3851), .CLK(clk_in), .RSTB(n7146), .Q(
        \FIFO[22][24] ) );
  DFFARX1 \FIFO_reg[22][23]  ( .D(n3850), .CLK(clk_in), .RSTB(n7146), .Q(
        \FIFO[22][23] ) );
  DFFARX1 \FIFO_reg[22][22]  ( .D(n3849), .CLK(clk_in), .RSTB(n7146), .Q(
        \FIFO[22][22] ) );
  DFFARX1 \FIFO_reg[22][21]  ( .D(n3848), .CLK(clk_in), .RSTB(n7146), .Q(
        \FIFO[22][21] ) );
  DFFARX1 \FIFO_reg[22][20]  ( .D(n3847), .CLK(clk_in), .RSTB(n7146), .Q(
        \FIFO[22][20] ) );
  DFFARX1 \FIFO_reg[22][19]  ( .D(n3846), .CLK(clk_in), .RSTB(n7146), .Q(
        \FIFO[22][19] ) );
  DFFARX1 \FIFO_reg[22][18]  ( .D(n3845), .CLK(clk_in), .RSTB(n7146), .Q(
        \FIFO[22][18] ) );
  DFFARX1 \FIFO_reg[22][17]  ( .D(n3844), .CLK(clk_in), .RSTB(n7146), .Q(
        \FIFO[22][17] ) );
  DFFARX1 \FIFO_reg[22][16]  ( .D(n3843), .CLK(clk_in), .RSTB(n7146), .Q(
        \FIFO[22][16] ) );
  DFFARX1 \FIFO_reg[22][15]  ( .D(n3842), .CLK(clk_in), .RSTB(n7146), .Q(
        \FIFO[22][15] ) );
  DFFARX1 \FIFO_reg[22][14]  ( .D(n3841), .CLK(clk_in), .RSTB(n7146), .Q(
        \FIFO[22][14] ) );
  DFFARX1 \FIFO_reg[22][13]  ( .D(n3840), .CLK(clk_in), .RSTB(n7146), .Q(
        \FIFO[22][13] ) );
  DFFARX1 \FIFO_reg[22][12]  ( .D(n3839), .CLK(clk_in), .RSTB(n7146), .Q(
        \FIFO[22][12] ) );
  DFFARX1 \FIFO_reg[22][11]  ( .D(n3838), .CLK(clk_in), .RSTB(n7146), .Q(
        \FIFO[22][11] ) );
  DFFARX1 \FIFO_reg[22][10]  ( .D(n3837), .CLK(clk_in), .RSTB(n7146), .Q(
        \FIFO[22][10] ) );
  DFFARX1 \FIFO_reg[22][9]  ( .D(n3836), .CLK(clk_in), .RSTB(n7147), .Q(
        \FIFO[22][9] ) );
  DFFARX1 \FIFO_reg[22][8]  ( .D(n3835), .CLK(clk_in), .RSTB(n7147), .Q(
        \FIFO[22][8] ) );
  DFFARX1 \FIFO_reg[22][7]  ( .D(n3834), .CLK(clk_in), .RSTB(n7147), .Q(
        \FIFO[22][7] ) );
  DFFARX1 \FIFO_reg[22][6]  ( .D(n3833), .CLK(clk_in), .RSTB(n7147), .Q(
        \FIFO[22][6] ) );
  DFFARX1 \FIFO_reg[22][5]  ( .D(n3832), .CLK(clk_in), .RSTB(n7147), .Q(
        \FIFO[22][5] ) );
  DFFARX1 \FIFO_reg[22][4]  ( .D(n3831), .CLK(clk_in), .RSTB(n7147), .Q(
        \FIFO[22][4] ) );
  DFFARX1 \FIFO_reg[22][3]  ( .D(n3830), .CLK(clk_in), .RSTB(n7147), .Q(
        \FIFO[22][3] ) );
  DFFARX1 \FIFO_reg[22][2]  ( .D(n3829), .CLK(clk_in), .RSTB(n7147), .Q(
        \FIFO[22][2] ) );
  DFFARX1 \FIFO_reg[22][1]  ( .D(n3828), .CLK(clk_in), .RSTB(n7147), .Q(
        \FIFO[22][1] ) );
  DFFARX1 \FIFO_reg[22][0]  ( .D(n3827), .CLK(clk_in), .RSTB(n7147), .Q(
        \FIFO[22][0] ) );
  DFFARX1 \FIFO_reg[23][31]  ( .D(n3826), .CLK(clk_in), .RSTB(n7147), .Q(
        \FIFO[23][31] ) );
  DFFARX1 \FIFO_reg[23][30]  ( .D(n3825), .CLK(clk_in), .RSTB(n7147), .Q(
        \FIFO[23][30] ) );
  DFFARX1 \FIFO_reg[23][29]  ( .D(n3824), .CLK(clk_in), .RSTB(n7147), .Q(
        \FIFO[23][29] ) );
  DFFARX1 \FIFO_reg[23][28]  ( .D(n3823), .CLK(clk_in), .RSTB(n7147), .Q(
        \FIFO[23][28] ) );
  DFFARX1 \FIFO_reg[23][27]  ( .D(n3822), .CLK(clk_in), .RSTB(n7147), .Q(
        \FIFO[23][27] ) );
  DFFARX1 \FIFO_reg[23][26]  ( .D(n3821), .CLK(clk_in), .RSTB(n7147), .Q(
        \FIFO[23][26] ) );
  DFFARX1 \FIFO_reg[23][25]  ( .D(n3820), .CLK(clk_in), .RSTB(n7147), .Q(
        \FIFO[23][25] ) );
  DFFARX1 \FIFO_reg[23][24]  ( .D(n3819), .CLK(clk_in), .RSTB(n7147), .Q(
        \FIFO[23][24] ) );
  DFFARX1 \FIFO_reg[23][23]  ( .D(n3818), .CLK(clk_in), .RSTB(n7148), .Q(
        \FIFO[23][23] ) );
  DFFARX1 \FIFO_reg[23][22]  ( .D(n3817), .CLK(clk_in), .RSTB(n7148), .Q(
        \FIFO[23][22] ) );
  DFFARX1 \FIFO_reg[23][21]  ( .D(n3816), .CLK(clk_in), .RSTB(n7148), .Q(
        \FIFO[23][21] ) );
  DFFARX1 \FIFO_reg[23][20]  ( .D(n3815), .CLK(clk_in), .RSTB(n7148), .Q(
        \FIFO[23][20] ) );
  DFFARX1 \FIFO_reg[23][19]  ( .D(n3814), .CLK(clk_in), .RSTB(n7148), .Q(
        \FIFO[23][19] ) );
  DFFARX1 \FIFO_reg[23][18]  ( .D(n3813), .CLK(clk_in), .RSTB(n7148), .Q(
        \FIFO[23][18] ) );
  DFFARX1 \FIFO_reg[23][17]  ( .D(n3812), .CLK(clk_in), .RSTB(n7148), .Q(
        \FIFO[23][17] ) );
  DFFARX1 \FIFO_reg[23][16]  ( .D(n3811), .CLK(clk_in), .RSTB(n7148), .Q(
        \FIFO[23][16] ) );
  DFFARX1 \FIFO_reg[23][15]  ( .D(n3810), .CLK(clk_in), .RSTB(n7148), .Q(
        \FIFO[23][15] ) );
  DFFARX1 \FIFO_reg[23][14]  ( .D(n3809), .CLK(clk_in), .RSTB(n7148), .Q(
        \FIFO[23][14] ) );
  DFFARX1 \FIFO_reg[23][13]  ( .D(n3808), .CLK(clk_in), .RSTB(n7148), .Q(
        \FIFO[23][13] ) );
  DFFARX1 \FIFO_reg[23][12]  ( .D(n3807), .CLK(clk_in), .RSTB(n7148), .Q(
        \FIFO[23][12] ) );
  DFFARX1 \FIFO_reg[23][11]  ( .D(n3806), .CLK(clk_in), .RSTB(n7148), .Q(
        \FIFO[23][11] ) );
  DFFARX1 \FIFO_reg[23][10]  ( .D(n3805), .CLK(clk_in), .RSTB(n7148), .Q(
        \FIFO[23][10] ) );
  DFFARX1 \FIFO_reg[23][9]  ( .D(n3804), .CLK(clk_in), .RSTB(n7148), .Q(
        \FIFO[23][9] ) );
  DFFARX1 \FIFO_reg[23][8]  ( .D(n3803), .CLK(clk_in), .RSTB(n7148), .Q(
        \FIFO[23][8] ) );
  DFFARX1 \FIFO_reg[23][7]  ( .D(n3802), .CLK(clk_in), .RSTB(n7148), .Q(
        \FIFO[23][7] ) );
  DFFARX1 \FIFO_reg[23][6]  ( .D(n3801), .CLK(clk_in), .RSTB(n7148), .Q(
        \FIFO[23][6] ) );
  DFFARX1 \FIFO_reg[23][5]  ( .D(n3800), .CLK(clk_in), .RSTB(n7149), .Q(
        \FIFO[23][5] ) );
  DFFARX1 \FIFO_reg[23][4]  ( .D(n3799), .CLK(clk_in), .RSTB(n7149), .Q(
        \FIFO[23][4] ) );
  DFFARX1 \FIFO_reg[23][3]  ( .D(n3798), .CLK(clk_in), .RSTB(n7149), .Q(
        \FIFO[23][3] ) );
  DFFARX1 \FIFO_reg[23][2]  ( .D(n3797), .CLK(clk_in), .RSTB(n7149), .Q(
        \FIFO[23][2] ) );
  DFFARX1 \FIFO_reg[23][1]  ( .D(n3796), .CLK(clk_in), .RSTB(n7149), .Q(
        \FIFO[23][1] ) );
  DFFARX1 \FIFO_reg[23][0]  ( .D(n3795), .CLK(clk_in), .RSTB(n7149), .Q(
        \FIFO[23][0] ) );
  DFFARX1 \FIFO_reg[24][31]  ( .D(n3794), .CLK(clk_in), .RSTB(n7149), .Q(
        \FIFO[24][31] ) );
  DFFARX1 \FIFO_reg[24][30]  ( .D(n3793), .CLK(clk_in), .RSTB(n7149), .Q(
        \FIFO[24][30] ) );
  DFFARX1 \FIFO_reg[24][29]  ( .D(n3792), .CLK(clk_in), .RSTB(n7149), .Q(
        \FIFO[24][29] ) );
  DFFARX1 \FIFO_reg[24][28]  ( .D(n3791), .CLK(clk_in), .RSTB(n7149), .Q(
        \FIFO[24][28] ) );
  DFFARX1 \FIFO_reg[24][27]  ( .D(n3790), .CLK(clk_in), .RSTB(n7149), .Q(
        \FIFO[24][27] ) );
  DFFARX1 \FIFO_reg[24][26]  ( .D(n3789), .CLK(clk_in), .RSTB(n7149), .Q(
        \FIFO[24][26] ) );
  DFFARX1 \FIFO_reg[24][25]  ( .D(n3788), .CLK(clk_in), .RSTB(n7149), .Q(
        \FIFO[24][25] ) );
  DFFARX1 \FIFO_reg[24][24]  ( .D(n3787), .CLK(clk_in), .RSTB(n7149), .Q(
        \FIFO[24][24] ) );
  DFFARX1 \FIFO_reg[24][23]  ( .D(n3786), .CLK(clk_in), .RSTB(n7149), .Q(
        \FIFO[24][23] ) );
  DFFARX1 \FIFO_reg[24][22]  ( .D(n3785), .CLK(clk_in), .RSTB(n7149), .Q(
        \FIFO[24][22] ) );
  DFFARX1 \FIFO_reg[24][21]  ( .D(n3784), .CLK(clk_in), .RSTB(n7149), .Q(
        \FIFO[24][21] ) );
  DFFARX1 \FIFO_reg[24][20]  ( .D(n3783), .CLK(clk_in), .RSTB(n7149), .Q(
        \FIFO[24][20] ) );
  DFFARX1 \FIFO_reg[24][19]  ( .D(n3782), .CLK(clk_in), .RSTB(n7150), .Q(
        \FIFO[24][19] ) );
  DFFARX1 \FIFO_reg[24][18]  ( .D(n3781), .CLK(clk_in), .RSTB(n7150), .Q(
        \FIFO[24][18] ) );
  DFFARX1 \FIFO_reg[24][17]  ( .D(n3780), .CLK(clk_in), .RSTB(n7150), .Q(
        \FIFO[24][17] ) );
  DFFARX1 \FIFO_reg[24][16]  ( .D(n3779), .CLK(clk_in), .RSTB(n7150), .Q(
        \FIFO[24][16] ) );
  DFFARX1 \FIFO_reg[24][15]  ( .D(n3778), .CLK(clk_in), .RSTB(n7150), .Q(
        \FIFO[24][15] ) );
  DFFARX1 \FIFO_reg[24][14]  ( .D(n3777), .CLK(clk_in), .RSTB(n7150), .Q(
        \FIFO[24][14] ) );
  DFFARX1 \FIFO_reg[24][13]  ( .D(n3776), .CLK(clk_in), .RSTB(n7150), .Q(
        \FIFO[24][13] ) );
  DFFARX1 \FIFO_reg[24][12]  ( .D(n3775), .CLK(clk_in), .RSTB(n7150), .Q(
        \FIFO[24][12] ) );
  DFFARX1 \FIFO_reg[24][11]  ( .D(n3774), .CLK(clk_in), .RSTB(n7150), .Q(
        \FIFO[24][11] ) );
  DFFARX1 \FIFO_reg[24][10]  ( .D(n3773), .CLK(clk_in), .RSTB(n7150), .Q(
        \FIFO[24][10] ) );
  DFFARX1 \FIFO_reg[24][9]  ( .D(n3772), .CLK(clk_in), .RSTB(n7150), .Q(
        \FIFO[24][9] ) );
  DFFARX1 \FIFO_reg[24][8]  ( .D(n3771), .CLK(clk_in), .RSTB(n7150), .Q(
        \FIFO[24][8] ) );
  DFFARX1 \FIFO_reg[24][7]  ( .D(n3770), .CLK(clk_in), .RSTB(n7150), .Q(
        \FIFO[24][7] ) );
  DFFARX1 \FIFO_reg[24][6]  ( .D(n3769), .CLK(clk_in), .RSTB(n7150), .Q(
        \FIFO[24][6] ) );
  DFFARX1 \FIFO_reg[24][5]  ( .D(n3768), .CLK(clk_in), .RSTB(n7150), .Q(
        \FIFO[24][5] ) );
  DFFARX1 \FIFO_reg[24][4]  ( .D(n3767), .CLK(clk_in), .RSTB(n7150), .Q(
        \FIFO[24][4] ) );
  DFFARX1 \FIFO_reg[24][3]  ( .D(n3766), .CLK(clk_in), .RSTB(n7150), .Q(
        \FIFO[24][3] ) );
  DFFARX1 \FIFO_reg[24][2]  ( .D(n3765), .CLK(clk_in), .RSTB(n7150), .Q(
        \FIFO[24][2] ) );
  DFFARX1 \FIFO_reg[24][1]  ( .D(n3764), .CLK(clk_in), .RSTB(n7151), .Q(
        \FIFO[24][1] ) );
  DFFARX1 \FIFO_reg[24][0]  ( .D(n3763), .CLK(clk_in), .RSTB(n7151), .Q(
        \FIFO[24][0] ) );
  DFFARX1 \FIFO_reg[25][31]  ( .D(n3762), .CLK(clk_in), .RSTB(n7151), .Q(
        \FIFO[25][31] ) );
  DFFARX1 \FIFO_reg[25][30]  ( .D(n3761), .CLK(clk_in), .RSTB(n7151), .Q(
        \FIFO[25][30] ) );
  DFFARX1 \FIFO_reg[25][29]  ( .D(n3760), .CLK(clk_in), .RSTB(n7151), .Q(
        \FIFO[25][29] ) );
  DFFARX1 \FIFO_reg[25][28]  ( .D(n3759), .CLK(clk_in), .RSTB(n7151), .Q(
        \FIFO[25][28] ) );
  DFFARX1 \FIFO_reg[25][27]  ( .D(n3758), .CLK(clk_in), .RSTB(n7151), .Q(
        \FIFO[25][27] ) );
  DFFARX1 \FIFO_reg[25][26]  ( .D(n3757), .CLK(clk_in), .RSTB(n7151), .Q(
        \FIFO[25][26] ) );
  DFFARX1 \FIFO_reg[25][25]  ( .D(n3756), .CLK(clk_in), .RSTB(n7151), .Q(
        \FIFO[25][25] ) );
  DFFARX1 \FIFO_reg[25][24]  ( .D(n3755), .CLK(clk_in), .RSTB(n7151), .Q(
        \FIFO[25][24] ) );
  DFFARX1 \FIFO_reg[25][23]  ( .D(n3754), .CLK(clk_in), .RSTB(n7151), .Q(
        \FIFO[25][23] ) );
  DFFARX1 \FIFO_reg[25][22]  ( .D(n3753), .CLK(clk_in), .RSTB(n7151), .Q(
        \FIFO[25][22] ) );
  DFFARX1 \FIFO_reg[25][21]  ( .D(n3752), .CLK(clk_in), .RSTB(n7151), .Q(
        \FIFO[25][21] ) );
  DFFARX1 \FIFO_reg[25][20]  ( .D(n3751), .CLK(clk_in), .RSTB(n7151), .Q(
        \FIFO[25][20] ) );
  DFFARX1 \FIFO_reg[25][19]  ( .D(n3750), .CLK(clk_in), .RSTB(n7151), .Q(
        \FIFO[25][19] ) );
  DFFARX1 \FIFO_reg[25][18]  ( .D(n3749), .CLK(clk_in), .RSTB(n7151), .Q(
        \FIFO[25][18] ) );
  DFFARX1 \FIFO_reg[25][17]  ( .D(n3748), .CLK(clk_in), .RSTB(n7151), .Q(
        \FIFO[25][17] ) );
  DFFARX1 \FIFO_reg[25][16]  ( .D(n3747), .CLK(clk_in), .RSTB(n7151), .Q(
        \FIFO[25][16] ) );
  DFFARX1 \FIFO_reg[25][15]  ( .D(n3746), .CLK(clk_in), .RSTB(n7152), .Q(
        \FIFO[25][15] ) );
  DFFARX1 \FIFO_reg[25][14]  ( .D(n3745), .CLK(clk_in), .RSTB(n7152), .Q(
        \FIFO[25][14] ) );
  DFFARX1 \FIFO_reg[25][13]  ( .D(n3744), .CLK(clk_in), .RSTB(n7152), .Q(
        \FIFO[25][13] ) );
  DFFARX1 \FIFO_reg[25][12]  ( .D(n3743), .CLK(clk_in), .RSTB(n7152), .Q(
        \FIFO[25][12] ) );
  DFFARX1 \FIFO_reg[25][11]  ( .D(n3742), .CLK(clk_in), .RSTB(n7152), .Q(
        \FIFO[25][11] ) );
  DFFARX1 \FIFO_reg[25][10]  ( .D(n3741), .CLK(clk_in), .RSTB(n7152), .Q(
        \FIFO[25][10] ) );
  DFFARX1 \FIFO_reg[25][9]  ( .D(n3740), .CLK(clk_in), .RSTB(n7152), .Q(
        \FIFO[25][9] ) );
  DFFARX1 \FIFO_reg[25][8]  ( .D(n3739), .CLK(clk_in), .RSTB(n7152), .Q(
        \FIFO[25][8] ) );
  DFFARX1 \FIFO_reg[25][7]  ( .D(n3738), .CLK(clk_in), .RSTB(n7152), .Q(
        \FIFO[25][7] ) );
  DFFARX1 \FIFO_reg[25][6]  ( .D(n3737), .CLK(clk_in), .RSTB(n7152), .Q(
        \FIFO[25][6] ) );
  DFFARX1 \FIFO_reg[25][5]  ( .D(n3736), .CLK(clk_in), .RSTB(n7152), .Q(
        \FIFO[25][5] ) );
  DFFARX1 \FIFO_reg[25][4]  ( .D(n3735), .CLK(clk_in), .RSTB(n7152), .Q(
        \FIFO[25][4] ) );
  DFFARX1 \FIFO_reg[25][3]  ( .D(n3734), .CLK(clk_in), .RSTB(n7152), .Q(
        \FIFO[25][3] ) );
  DFFARX1 \FIFO_reg[25][2]  ( .D(n3733), .CLK(clk_in), .RSTB(n7152), .Q(
        \FIFO[25][2] ) );
  DFFARX1 \FIFO_reg[25][1]  ( .D(n3732), .CLK(clk_in), .RSTB(n7152), .Q(
        \FIFO[25][1] ) );
  DFFARX1 \FIFO_reg[25][0]  ( .D(n3731), .CLK(clk_in), .RSTB(n7152), .Q(
        \FIFO[25][0] ) );
  DFFARX1 \FIFO_reg[26][31]  ( .D(n3730), .CLK(clk_in), .RSTB(n7152), .Q(
        \FIFO[26][31] ) );
  DFFARX1 \FIFO_reg[26][30]  ( .D(n3729), .CLK(clk_in), .RSTB(n7152), .Q(
        \FIFO[26][30] ) );
  DFFARX1 \FIFO_reg[26][29]  ( .D(n3728), .CLK(clk_in), .RSTB(n7153), .Q(
        \FIFO[26][29] ) );
  DFFARX1 \FIFO_reg[26][28]  ( .D(n3727), .CLK(clk_in), .RSTB(n7153), .Q(
        \FIFO[26][28] ) );
  DFFARX1 \FIFO_reg[26][27]  ( .D(n3726), .CLK(clk_in), .RSTB(n7153), .Q(
        \FIFO[26][27] ) );
  DFFARX1 \FIFO_reg[26][26]  ( .D(n3725), .CLK(clk_in), .RSTB(n7153), .Q(
        \FIFO[26][26] ) );
  DFFARX1 \FIFO_reg[26][25]  ( .D(n3724), .CLK(clk_in), .RSTB(n7153), .Q(
        \FIFO[26][25] ) );
  DFFARX1 \FIFO_reg[26][24]  ( .D(n3723), .CLK(clk_in), .RSTB(n7153), .Q(
        \FIFO[26][24] ) );
  DFFARX1 \FIFO_reg[26][23]  ( .D(n3722), .CLK(clk_in), .RSTB(n7153), .Q(
        \FIFO[26][23] ) );
  DFFARX1 \FIFO_reg[26][22]  ( .D(n3721), .CLK(clk_in), .RSTB(n7153), .Q(
        \FIFO[26][22] ) );
  DFFARX1 \FIFO_reg[26][21]  ( .D(n3720), .CLK(clk_in), .RSTB(n7153), .Q(
        \FIFO[26][21] ) );
  DFFARX1 \FIFO_reg[26][20]  ( .D(n3719), .CLK(clk_in), .RSTB(n7153), .Q(
        \FIFO[26][20] ) );
  DFFARX1 \FIFO_reg[26][19]  ( .D(n3718), .CLK(clk_in), .RSTB(n7153), .Q(
        \FIFO[26][19] ) );
  DFFARX1 \FIFO_reg[26][18]  ( .D(n3717), .CLK(clk_in), .RSTB(n7153), .Q(
        \FIFO[26][18] ) );
  DFFARX1 \FIFO_reg[26][17]  ( .D(n3716), .CLK(clk_in), .RSTB(n7153), .Q(
        \FIFO[26][17] ) );
  DFFARX1 \FIFO_reg[26][16]  ( .D(n3715), .CLK(clk_in), .RSTB(n7153), .Q(
        \FIFO[26][16] ) );
  DFFARX1 \FIFO_reg[26][15]  ( .D(n3714), .CLK(clk_in), .RSTB(n7153), .Q(
        \FIFO[26][15] ) );
  DFFARX1 \FIFO_reg[26][14]  ( .D(n3713), .CLK(clk_in), .RSTB(n7153), .Q(
        \FIFO[26][14] ) );
  DFFARX1 \FIFO_reg[26][13]  ( .D(n3712), .CLK(clk_in), .RSTB(n7153), .Q(
        \FIFO[26][13] ) );
  DFFARX1 \FIFO_reg[26][12]  ( .D(n3711), .CLK(clk_in), .RSTB(n7153), .Q(
        \FIFO[26][12] ) );
  DFFARX1 \FIFO_reg[26][11]  ( .D(n3710), .CLK(clk_in), .RSTB(n7154), .Q(
        \FIFO[26][11] ) );
  DFFARX1 \FIFO_reg[26][10]  ( .D(n3709), .CLK(clk_in), .RSTB(n7154), .Q(
        \FIFO[26][10] ) );
  DFFARX1 \FIFO_reg[26][9]  ( .D(n3708), .CLK(clk_in), .RSTB(n7154), .Q(
        \FIFO[26][9] ) );
  DFFARX1 \FIFO_reg[26][8]  ( .D(n3707), .CLK(clk_in), .RSTB(n7154), .Q(
        \FIFO[26][8] ) );
  DFFARX1 \FIFO_reg[26][7]  ( .D(n3706), .CLK(clk_in), .RSTB(n7154), .Q(
        \FIFO[26][7] ) );
  DFFARX1 \FIFO_reg[26][6]  ( .D(n3705), .CLK(clk_in), .RSTB(n7154), .Q(
        \FIFO[26][6] ) );
  DFFARX1 \FIFO_reg[26][5]  ( .D(n3704), .CLK(clk_in), .RSTB(n7154), .Q(
        \FIFO[26][5] ) );
  DFFARX1 \FIFO_reg[26][4]  ( .D(n3703), .CLK(clk_in), .RSTB(n7154), .Q(
        \FIFO[26][4] ) );
  DFFARX1 \FIFO_reg[26][3]  ( .D(n3702), .CLK(clk_in), .RSTB(n7154), .Q(
        \FIFO[26][3] ) );
  DFFARX1 \FIFO_reg[26][2]  ( .D(n3701), .CLK(clk_in), .RSTB(n7154), .Q(
        \FIFO[26][2] ) );
  DFFARX1 \FIFO_reg[26][1]  ( .D(n3700), .CLK(clk_in), .RSTB(n7154), .Q(
        \FIFO[26][1] ) );
  DFFARX1 \FIFO_reg[26][0]  ( .D(n3699), .CLK(clk_in), .RSTB(n7154), .Q(
        \FIFO[26][0] ) );
  DFFARX1 \FIFO_reg[27][31]  ( .D(n3698), .CLK(clk_in), .RSTB(n7154), .Q(
        \FIFO[27][31] ) );
  DFFARX1 \FIFO_reg[27][30]  ( .D(n3697), .CLK(clk_in), .RSTB(n7154), .Q(
        \FIFO[27][30] ) );
  DFFARX1 \FIFO_reg[27][29]  ( .D(n3696), .CLK(clk_in), .RSTB(n7154), .Q(
        \FIFO[27][29] ) );
  DFFARX1 \FIFO_reg[27][28]  ( .D(n3695), .CLK(clk_in), .RSTB(n7154), .Q(
        \FIFO[27][28] ) );
  DFFARX1 \FIFO_reg[27][27]  ( .D(n3694), .CLK(clk_in), .RSTB(n7154), .Q(
        \FIFO[27][27] ) );
  DFFARX1 \FIFO_reg[27][26]  ( .D(n3693), .CLK(clk_in), .RSTB(n7154), .Q(
        \FIFO[27][26] ) );
  DFFARX1 \FIFO_reg[27][25]  ( .D(n3692), .CLK(clk_in), .RSTB(n7155), .Q(
        \FIFO[27][25] ) );
  DFFARX1 \FIFO_reg[27][24]  ( .D(n3691), .CLK(clk_in), .RSTB(n7155), .Q(
        \FIFO[27][24] ) );
  DFFARX1 \FIFO_reg[27][23]  ( .D(n3690), .CLK(clk_in), .RSTB(n7155), .Q(
        \FIFO[27][23] ) );
  DFFARX1 \FIFO_reg[27][22]  ( .D(n3689), .CLK(clk_in), .RSTB(n7155), .Q(
        \FIFO[27][22] ) );
  DFFARX1 \FIFO_reg[27][21]  ( .D(n3688), .CLK(clk_in), .RSTB(n7155), .Q(
        \FIFO[27][21] ) );
  DFFARX1 \FIFO_reg[27][20]  ( .D(n3687), .CLK(clk_in), .RSTB(n7155), .Q(
        \FIFO[27][20] ) );
  DFFARX1 \FIFO_reg[27][19]  ( .D(n3686), .CLK(clk_in), .RSTB(n7155), .Q(
        \FIFO[27][19] ) );
  DFFARX1 \FIFO_reg[27][18]  ( .D(n3685), .CLK(clk_in), .RSTB(n7155), .Q(
        \FIFO[27][18] ) );
  DFFARX1 \FIFO_reg[27][17]  ( .D(n3684), .CLK(clk_in), .RSTB(n7155), .Q(
        \FIFO[27][17] ) );
  DFFARX1 \FIFO_reg[27][16]  ( .D(n3683), .CLK(clk_in), .RSTB(n7155), .Q(
        \FIFO[27][16] ) );
  DFFARX1 \FIFO_reg[27][15]  ( .D(n3682), .CLK(clk_in), .RSTB(n7155), .Q(
        \FIFO[27][15] ) );
  DFFARX1 \FIFO_reg[27][14]  ( .D(n3681), .CLK(clk_in), .RSTB(n7155), .Q(
        \FIFO[27][14] ) );
  DFFARX1 \FIFO_reg[27][13]  ( .D(n3680), .CLK(clk_in), .RSTB(n7155), .Q(
        \FIFO[27][13] ) );
  DFFARX1 \FIFO_reg[27][12]  ( .D(n3679), .CLK(clk_in), .RSTB(n7155), .Q(
        \FIFO[27][12] ) );
  DFFARX1 \FIFO_reg[27][11]  ( .D(n3678), .CLK(clk_in), .RSTB(n7155), .Q(
        \FIFO[27][11] ) );
  DFFARX1 \FIFO_reg[27][10]  ( .D(n3677), .CLK(clk_in), .RSTB(n7155), .Q(
        \FIFO[27][10] ) );
  DFFARX1 \FIFO_reg[27][9]  ( .D(n3676), .CLK(clk_in), .RSTB(n7155), .Q(
        \FIFO[27][9] ) );
  DFFARX1 \FIFO_reg[27][8]  ( .D(n3675), .CLK(clk_in), .RSTB(n7155), .Q(
        \FIFO[27][8] ) );
  DFFARX1 \FIFO_reg[27][7]  ( .D(n3674), .CLK(clk_in), .RSTB(n7156), .Q(
        \FIFO[27][7] ) );
  DFFARX1 \FIFO_reg[27][6]  ( .D(n3673), .CLK(clk_in), .RSTB(n7156), .Q(
        \FIFO[27][6] ) );
  DFFARX1 \FIFO_reg[27][5]  ( .D(n3672), .CLK(clk_in), .RSTB(n7156), .Q(
        \FIFO[27][5] ) );
  DFFARX1 \FIFO_reg[27][4]  ( .D(n3671), .CLK(clk_in), .RSTB(n7156), .Q(
        \FIFO[27][4] ) );
  DFFARX1 \FIFO_reg[27][3]  ( .D(n3670), .CLK(clk_in), .RSTB(n7156), .Q(
        \FIFO[27][3] ) );
  DFFARX1 \FIFO_reg[27][2]  ( .D(n3669), .CLK(clk_in), .RSTB(n7156), .Q(
        \FIFO[27][2] ) );
  DFFARX1 \FIFO_reg[27][1]  ( .D(n3668), .CLK(clk_in), .RSTB(n7156), .Q(
        \FIFO[27][1] ) );
  DFFARX1 \FIFO_reg[27][0]  ( .D(n3667), .CLK(clk_in), .RSTB(n7156), .Q(
        \FIFO[27][0] ) );
  DFFARX1 \FIFO_reg[28][31]  ( .D(n3666), .CLK(clk_in), .RSTB(n7156), .Q(
        \FIFO[28][31] ) );
  DFFARX1 \FIFO_reg[28][30]  ( .D(n3665), .CLK(clk_in), .RSTB(n7156), .Q(
        \FIFO[28][30] ) );
  DFFARX1 \FIFO_reg[28][29]  ( .D(n3664), .CLK(clk_in), .RSTB(n7156), .Q(
        \FIFO[28][29] ) );
  DFFARX1 \FIFO_reg[28][28]  ( .D(n3663), .CLK(clk_in), .RSTB(n7156), .Q(
        \FIFO[28][28] ) );
  DFFARX1 \FIFO_reg[28][27]  ( .D(n3662), .CLK(clk_in), .RSTB(n7156), .Q(
        \FIFO[28][27] ) );
  DFFARX1 \FIFO_reg[28][26]  ( .D(n3661), .CLK(clk_in), .RSTB(n7156), .Q(
        \FIFO[28][26] ) );
  DFFARX1 \FIFO_reg[28][25]  ( .D(n3660), .CLK(clk_in), .RSTB(n7156), .Q(
        \FIFO[28][25] ) );
  DFFARX1 \FIFO_reg[28][24]  ( .D(n3659), .CLK(clk_in), .RSTB(n7156), .Q(
        \FIFO[28][24] ) );
  DFFARX1 \FIFO_reg[28][23]  ( .D(n3658), .CLK(clk_in), .RSTB(n7156), .Q(
        \FIFO[28][23] ) );
  DFFARX1 \FIFO_reg[28][22]  ( .D(n3657), .CLK(clk_in), .RSTB(n7156), .Q(
        \FIFO[28][22] ) );
  DFFARX1 \FIFO_reg[28][21]  ( .D(n3656), .CLK(clk_in), .RSTB(n7157), .Q(
        \FIFO[28][21] ) );
  DFFARX1 \FIFO_reg[28][20]  ( .D(n3655), .CLK(clk_in), .RSTB(n7157), .Q(
        \FIFO[28][20] ) );
  DFFARX1 \FIFO_reg[28][19]  ( .D(n3654), .CLK(clk_in), .RSTB(n7157), .Q(
        \FIFO[28][19] ) );
  DFFARX1 \FIFO_reg[28][18]  ( .D(n3653), .CLK(clk_in), .RSTB(n7157), .Q(
        \FIFO[28][18] ) );
  DFFARX1 \FIFO_reg[28][17]  ( .D(n3652), .CLK(clk_in), .RSTB(n7157), .Q(
        \FIFO[28][17] ) );
  DFFARX1 \FIFO_reg[28][16]  ( .D(n3651), .CLK(clk_in), .RSTB(n7157), .Q(
        \FIFO[28][16] ) );
  DFFARX1 \FIFO_reg[28][15]  ( .D(n3650), .CLK(clk_in), .RSTB(n7157), .Q(
        \FIFO[28][15] ) );
  DFFARX1 \FIFO_reg[28][14]  ( .D(n3649), .CLK(clk_in), .RSTB(n7157), .Q(
        \FIFO[28][14] ) );
  DFFARX1 \FIFO_reg[28][13]  ( .D(n3648), .CLK(clk_in), .RSTB(n7157), .Q(
        \FIFO[28][13] ) );
  DFFARX1 \FIFO_reg[28][12]  ( .D(n3647), .CLK(clk_in), .RSTB(n7157), .Q(
        \FIFO[28][12] ) );
  DFFARX1 \FIFO_reg[28][11]  ( .D(n3646), .CLK(clk_in), .RSTB(n7157), .Q(
        \FIFO[28][11] ) );
  DFFARX1 \FIFO_reg[28][10]  ( .D(n3645), .CLK(clk_in), .RSTB(n7157), .Q(
        \FIFO[28][10] ) );
  DFFARX1 \FIFO_reg[28][9]  ( .D(n3644), .CLK(clk_in), .RSTB(n7157), .Q(
        \FIFO[28][9] ) );
  DFFARX1 \FIFO_reg[28][8]  ( .D(n3643), .CLK(clk_in), .RSTB(n7157), .Q(
        \FIFO[28][8] ) );
  DFFARX1 \FIFO_reg[28][7]  ( .D(n3642), .CLK(clk_in), .RSTB(n7157), .Q(
        \FIFO[28][7] ) );
  DFFARX1 \FIFO_reg[28][6]  ( .D(n3641), .CLK(clk_in), .RSTB(n7157), .Q(
        \FIFO[28][6] ) );
  DFFARX1 \FIFO_reg[28][5]  ( .D(n3640), .CLK(clk_in), .RSTB(n7157), .Q(
        \FIFO[28][5] ) );
  DFFARX1 \FIFO_reg[28][4]  ( .D(n3639), .CLK(clk_in), .RSTB(n7157), .Q(
        \FIFO[28][4] ) );
  DFFARX1 \FIFO_reg[28][3]  ( .D(n3638), .CLK(clk_in), .RSTB(n7158), .Q(
        \FIFO[28][3] ) );
  DFFARX1 \FIFO_reg[28][2]  ( .D(n3637), .CLK(clk_in), .RSTB(n7158), .Q(
        \FIFO[28][2] ) );
  DFFARX1 \FIFO_reg[28][1]  ( .D(n3636), .CLK(clk_in), .RSTB(n7158), .Q(
        \FIFO[28][1] ) );
  DFFARX1 \FIFO_reg[28][0]  ( .D(n3635), .CLK(clk_in), .RSTB(n7158), .Q(
        \FIFO[28][0] ) );
  DFFARX1 \FIFO_reg[29][31]  ( .D(n3634), .CLK(clk_in), .RSTB(n7158), .Q(
        \FIFO[29][31] ) );
  DFFARX1 \FIFO_reg[29][30]  ( .D(n3633), .CLK(clk_in), .RSTB(n7158), .Q(
        \FIFO[29][30] ) );
  DFFARX1 \FIFO_reg[29][29]  ( .D(n3632), .CLK(clk_in), .RSTB(n7158), .Q(
        \FIFO[29][29] ) );
  DFFARX1 \FIFO_reg[29][28]  ( .D(n3631), .CLK(clk_in), .RSTB(n7158), .Q(
        \FIFO[29][28] ) );
  DFFARX1 \FIFO_reg[29][27]  ( .D(n3630), .CLK(clk_in), .RSTB(n7158), .Q(
        \FIFO[29][27] ) );
  DFFARX1 \FIFO_reg[29][26]  ( .D(n3629), .CLK(clk_in), .RSTB(n7158), .Q(
        \FIFO[29][26] ) );
  DFFARX1 \FIFO_reg[29][25]  ( .D(n3628), .CLK(clk_in), .RSTB(n7158), .Q(
        \FIFO[29][25] ) );
  DFFARX1 \FIFO_reg[29][24]  ( .D(n3627), .CLK(clk_in), .RSTB(n7158), .Q(
        \FIFO[29][24] ) );
  DFFARX1 \FIFO_reg[29][23]  ( .D(n3626), .CLK(clk_in), .RSTB(n7158), .Q(
        \FIFO[29][23] ) );
  DFFARX1 \FIFO_reg[29][22]  ( .D(n3625), .CLK(clk_in), .RSTB(n7158), .Q(
        \FIFO[29][22] ) );
  DFFARX1 \FIFO_reg[29][21]  ( .D(n3624), .CLK(clk_in), .RSTB(n7158), .Q(
        \FIFO[29][21] ) );
  DFFARX1 \FIFO_reg[29][20]  ( .D(n3623), .CLK(clk_in), .RSTB(n7158), .Q(
        \FIFO[29][20] ) );
  DFFARX1 \FIFO_reg[29][19]  ( .D(n3622), .CLK(clk_in), .RSTB(n7158), .Q(
        \FIFO[29][19] ) );
  DFFARX1 \FIFO_reg[29][18]  ( .D(n3621), .CLK(clk_in), .RSTB(n7158), .Q(
        \FIFO[29][18] ) );
  DFFARX1 \FIFO_reg[29][17]  ( .D(n3620), .CLK(clk_in), .RSTB(n7159), .Q(
        \FIFO[29][17] ) );
  DFFARX1 \FIFO_reg[29][16]  ( .D(n3619), .CLK(clk_in), .RSTB(n7159), .Q(
        \FIFO[29][16] ) );
  DFFARX1 \FIFO_reg[29][15]  ( .D(n3618), .CLK(clk_in), .RSTB(n7159), .Q(
        \FIFO[29][15] ) );
  DFFARX1 \FIFO_reg[29][14]  ( .D(n3617), .CLK(clk_in), .RSTB(n7159), .Q(
        \FIFO[29][14] ) );
  DFFARX1 \FIFO_reg[29][13]  ( .D(n3616), .CLK(clk_in), .RSTB(n7159), .Q(
        \FIFO[29][13] ) );
  DFFARX1 \FIFO_reg[29][12]  ( .D(n3615), .CLK(clk_in), .RSTB(n7159), .Q(
        \FIFO[29][12] ) );
  DFFARX1 \FIFO_reg[29][11]  ( .D(n3614), .CLK(clk_in), .RSTB(n7159), .Q(
        \FIFO[29][11] ) );
  DFFARX1 \FIFO_reg[29][10]  ( .D(n3613), .CLK(clk_in), .RSTB(n7159), .Q(
        \FIFO[29][10] ) );
  DFFARX1 \FIFO_reg[29][9]  ( .D(n3612), .CLK(clk_in), .RSTB(n7159), .Q(
        \FIFO[29][9] ) );
  DFFARX1 \FIFO_reg[29][8]  ( .D(n3611), .CLK(clk_in), .RSTB(n7159), .Q(
        \FIFO[29][8] ) );
  DFFARX1 \FIFO_reg[29][7]  ( .D(n3610), .CLK(clk_in), .RSTB(n7159), .Q(
        \FIFO[29][7] ) );
  DFFARX1 \FIFO_reg[29][6]  ( .D(n3609), .CLK(clk_in), .RSTB(n7159), .Q(
        \FIFO[29][6] ) );
  DFFARX1 \FIFO_reg[29][5]  ( .D(n3608), .CLK(clk_in), .RSTB(n7159), .Q(
        \FIFO[29][5] ) );
  DFFARX1 \FIFO_reg[29][4]  ( .D(n3607), .CLK(clk_in), .RSTB(n7159), .Q(
        \FIFO[29][4] ) );
  DFFARX1 \FIFO_reg[29][3]  ( .D(n3606), .CLK(clk_in), .RSTB(n7159), .Q(
        \FIFO[29][3] ) );
  DFFARX1 \FIFO_reg[29][2]  ( .D(n3605), .CLK(clk_in), .RSTB(n7159), .Q(
        \FIFO[29][2] ) );
  DFFARX1 \FIFO_reg[29][1]  ( .D(n3604), .CLK(clk_in), .RSTB(n7159), .Q(
        \FIFO[29][1] ) );
  DFFARX1 \FIFO_reg[29][0]  ( .D(n3603), .CLK(clk_in), .RSTB(n7159), .Q(
        \FIFO[29][0] ) );
  DFFARX1 \FIFO_reg[30][31]  ( .D(n3602), .CLK(clk_in), .RSTB(n7160), .Q(
        \FIFO[30][31] ) );
  DFFARX1 \FIFO_reg[30][30]  ( .D(n3601), .CLK(clk_in), .RSTB(n7160), .Q(
        \FIFO[30][30] ) );
  DFFARX1 \FIFO_reg[30][29]  ( .D(n3600), .CLK(clk_in), .RSTB(n7160), .Q(
        \FIFO[30][29] ) );
  DFFARX1 \FIFO_reg[30][28]  ( .D(n3599), .CLK(clk_in), .RSTB(n7160), .Q(
        \FIFO[30][28] ) );
  DFFARX1 \FIFO_reg[30][27]  ( .D(n3598), .CLK(clk_in), .RSTB(n7160), .Q(
        \FIFO[30][27] ) );
  DFFARX1 \FIFO_reg[30][26]  ( .D(n3597), .CLK(clk_in), .RSTB(n7160), .Q(
        \FIFO[30][26] ) );
  DFFARX1 \FIFO_reg[30][25]  ( .D(n3596), .CLK(clk_in), .RSTB(n7160), .Q(
        \FIFO[30][25] ) );
  DFFARX1 \FIFO_reg[30][24]  ( .D(n3595), .CLK(clk_in), .RSTB(n7160), .Q(
        \FIFO[30][24] ) );
  DFFARX1 \FIFO_reg[30][23]  ( .D(n3594), .CLK(clk_in), .RSTB(n7160), .Q(
        \FIFO[30][23] ) );
  DFFARX1 \FIFO_reg[30][22]  ( .D(n3593), .CLK(clk_in), .RSTB(n7160), .Q(
        \FIFO[30][22] ) );
  DFFARX1 \FIFO_reg[30][21]  ( .D(n3592), .CLK(clk_in), .RSTB(n7160), .Q(
        \FIFO[30][21] ) );
  DFFARX1 \FIFO_reg[30][20]  ( .D(n3591), .CLK(clk_in), .RSTB(n7160), .Q(
        \FIFO[30][20] ) );
  DFFARX1 \FIFO_reg[30][19]  ( .D(n3590), .CLK(clk_in), .RSTB(n7160), .Q(
        \FIFO[30][19] ) );
  DFFARX1 \FIFO_reg[30][18]  ( .D(n3589), .CLK(clk_in), .RSTB(n7160), .Q(
        \FIFO[30][18] ) );
  DFFARX1 \FIFO_reg[30][17]  ( .D(n3588), .CLK(clk_in), .RSTB(n7160), .Q(
        \FIFO[30][17] ) );
  DFFARX1 \FIFO_reg[30][16]  ( .D(n3587), .CLK(clk_in), .RSTB(n7160), .Q(
        \FIFO[30][16] ) );
  DFFARX1 \FIFO_reg[30][15]  ( .D(n3586), .CLK(clk_in), .RSTB(n7160), .Q(
        \FIFO[30][15] ) );
  DFFARX1 \FIFO_reg[30][14]  ( .D(n3585), .CLK(clk_in), .RSTB(n7160), .Q(
        \FIFO[30][14] ) );
  DFFARX1 \FIFO_reg[30][13]  ( .D(n3584), .CLK(clk_in), .RSTB(n7161), .Q(
        \FIFO[30][13] ) );
  DFFARX1 \FIFO_reg[30][12]  ( .D(n3583), .CLK(clk_in), .RSTB(n7161), .Q(
        \FIFO[30][12] ) );
  DFFARX1 \FIFO_reg[30][11]  ( .D(n3582), .CLK(clk_in), .RSTB(n7161), .Q(
        \FIFO[30][11] ) );
  DFFARX1 \FIFO_reg[30][10]  ( .D(n3581), .CLK(clk_in), .RSTB(n7161), .Q(
        \FIFO[30][10] ) );
  DFFARX1 \FIFO_reg[30][9]  ( .D(n3580), .CLK(clk_in), .RSTB(n7161), .Q(
        \FIFO[30][9] ) );
  DFFARX1 \FIFO_reg[30][8]  ( .D(n3579), .CLK(clk_in), .RSTB(n7161), .Q(
        \FIFO[30][8] ) );
  DFFARX1 \FIFO_reg[30][7]  ( .D(n3578), .CLK(clk_in), .RSTB(n7161), .Q(
        \FIFO[30][7] ) );
  DFFARX1 \FIFO_reg[30][6]  ( .D(n3577), .CLK(clk_in), .RSTB(n7161), .Q(
        \FIFO[30][6] ) );
  DFFARX1 \FIFO_reg[30][5]  ( .D(n3576), .CLK(clk_in), .RSTB(n7161), .Q(
        \FIFO[30][5] ) );
  DFFARX1 \FIFO_reg[30][4]  ( .D(n3575), .CLK(clk_in), .RSTB(n7161), .Q(
        \FIFO[30][4] ) );
  DFFARX1 \FIFO_reg[30][3]  ( .D(n3574), .CLK(clk_in), .RSTB(n7161), .Q(
        \FIFO[30][3] ) );
  DFFARX1 \FIFO_reg[30][2]  ( .D(n3573), .CLK(clk_in), .RSTB(n7161), .Q(
        \FIFO[30][2] ) );
  DFFARX1 \FIFO_reg[30][1]  ( .D(n3572), .CLK(clk_in), .RSTB(n7161), .Q(
        \FIFO[30][1] ) );
  DFFARX1 \FIFO_reg[30][0]  ( .D(n3571), .CLK(clk_in), .RSTB(n7161), .Q(
        \FIFO[30][0] ) );
  DFFARX1 \FIFO_reg[31][31]  ( .D(n3570), .CLK(clk_in), .RSTB(n7161), .Q(
        \FIFO[31][31] ) );
  DFFARX1 \FIFO_reg[31][30]  ( .D(n3569), .CLK(clk_in), .RSTB(n7161), .Q(
        \FIFO[31][30] ) );
  DFFARX1 \FIFO_reg[31][29]  ( .D(n3568), .CLK(clk_in), .RSTB(n7161), .Q(
        \FIFO[31][29] ) );
  DFFARX1 \FIFO_reg[31][28]  ( .D(n3567), .CLK(clk_in), .RSTB(n7161), .Q(
        \FIFO[31][28] ) );
  DFFARX1 \FIFO_reg[31][27]  ( .D(n3566), .CLK(clk_in), .RSTB(n7162), .Q(
        \FIFO[31][27] ) );
  DFFARX1 \FIFO_reg[31][26]  ( .D(n3565), .CLK(clk_in), .RSTB(n7162), .Q(
        \FIFO[31][26] ) );
  DFFARX1 \FIFO_reg[31][25]  ( .D(n3564), .CLK(clk_in), .RSTB(n7162), .Q(
        \FIFO[31][25] ) );
  DFFARX1 \FIFO_reg[31][24]  ( .D(n3563), .CLK(clk_in), .RSTB(n7162), .Q(
        \FIFO[31][24] ) );
  DFFARX1 \FIFO_reg[31][23]  ( .D(n3562), .CLK(clk_in), .RSTB(n7162), .Q(
        \FIFO[31][23] ) );
  DFFARX1 \FIFO_reg[31][22]  ( .D(n3561), .CLK(clk_in), .RSTB(n7162), .Q(
        \FIFO[31][22] ) );
  DFFARX1 \FIFO_reg[31][21]  ( .D(n3560), .CLK(clk_in), .RSTB(n7162), .Q(
        \FIFO[31][21] ) );
  DFFARX1 \FIFO_reg[31][20]  ( .D(n3559), .CLK(clk_in), .RSTB(n7162), .Q(
        \FIFO[31][20] ) );
  DFFARX1 \FIFO_reg[31][19]  ( .D(n3558), .CLK(clk_in), .RSTB(n7162), .Q(
        \FIFO[31][19] ) );
  DFFARX1 \FIFO_reg[31][18]  ( .D(n3557), .CLK(clk_in), .RSTB(n7162), .Q(
        \FIFO[31][18] ) );
  DFFARX1 \FIFO_reg[31][17]  ( .D(n3556), .CLK(clk_in), .RSTB(n7162), .Q(
        \FIFO[31][17] ) );
  DFFARX1 \FIFO_reg[31][16]  ( .D(n3555), .CLK(clk_in), .RSTB(n7162), .Q(
        \FIFO[31][16] ) );
  DFFARX1 \FIFO_reg[31][15]  ( .D(n3554), .CLK(clk_in), .RSTB(n7162), .Q(
        \FIFO[31][15] ) );
  DFFARX1 \FIFO_reg[31][14]  ( .D(n3553), .CLK(clk_in), .RSTB(n7162), .Q(
        \FIFO[31][14] ) );
  DFFARX1 \FIFO_reg[31][13]  ( .D(n3552), .CLK(clk_in), .RSTB(n7162), .Q(
        \FIFO[31][13] ) );
  DFFARX1 \FIFO_reg[31][12]  ( .D(n3551), .CLK(clk_in), .RSTB(n7162), .Q(
        \FIFO[31][12] ) );
  DFFARX1 \FIFO_reg[31][11]  ( .D(n3550), .CLK(clk_in), .RSTB(n7162), .Q(
        \FIFO[31][11] ) );
  DFFARX1 \FIFO_reg[31][10]  ( .D(n3549), .CLK(clk_in), .RSTB(n7162), .Q(
        \FIFO[31][10] ) );
  DFFARX1 \FIFO_reg[31][9]  ( .D(n3548), .CLK(clk_in), .RSTB(n7163), .Q(
        \FIFO[31][9] ) );
  DFFARX1 \FIFO_reg[31][8]  ( .D(n3547), .CLK(clk_in), .RSTB(n7163), .Q(
        \FIFO[31][8] ) );
  DFFARX1 \FIFO_reg[31][7]  ( .D(n3546), .CLK(clk_in), .RSTB(n7163), .Q(
        \FIFO[31][7] ) );
  DFFARX1 \FIFO_reg[31][6]  ( .D(n3545), .CLK(clk_in), .RSTB(n7163), .Q(
        \FIFO[31][6] ) );
  DFFARX1 \FIFO_reg[31][5]  ( .D(n3544), .CLK(clk_in), .RSTB(n7163), .Q(
        \FIFO[31][5] ) );
  DFFARX1 \FIFO_reg[31][4]  ( .D(n3543), .CLK(clk_in), .RSTB(n7163), .Q(
        \FIFO[31][4] ) );
  DFFARX1 \FIFO_reg[31][3]  ( .D(n3542), .CLK(clk_in), .RSTB(n7163), .Q(
        \FIFO[31][3] ) );
  DFFARX1 \FIFO_reg[31][2]  ( .D(n3541), .CLK(clk_in), .RSTB(n7163), .Q(
        \FIFO[31][2] ) );
  DFFARX1 \FIFO_reg[31][1]  ( .D(n3540), .CLK(clk_in), .RSTB(n7163), .Q(
        \FIFO[31][1] ) );
  DFFARX1 \FIFO_reg[31][0]  ( .D(n3539), .CLK(clk_in), .RSTB(n7163), .Q(
        \FIFO[31][0] ) );
  DFFARX1 \FIFO_reg[32][31]  ( .D(n3538), .CLK(clk_in), .RSTB(n7163), .Q(
        \FIFO[32][31] ) );
  DFFARX1 \FIFO_reg[32][30]  ( .D(n3537), .CLK(clk_in), .RSTB(n7163), .Q(
        \FIFO[32][30] ) );
  DFFARX1 \FIFO_reg[32][29]  ( .D(n3536), .CLK(clk_in), .RSTB(n7163), .Q(
        \FIFO[32][29] ) );
  DFFARX1 \FIFO_reg[32][28]  ( .D(n3535), .CLK(clk_in), .RSTB(n7163), .Q(
        \FIFO[32][28] ) );
  DFFARX1 \FIFO_reg[32][27]  ( .D(n3534), .CLK(clk_in), .RSTB(n7163), .Q(
        \FIFO[32][27] ) );
  DFFARX1 \FIFO_reg[32][26]  ( .D(n3533), .CLK(clk_in), .RSTB(n7163), .Q(
        \FIFO[32][26] ) );
  DFFARX1 \FIFO_reg[32][25]  ( .D(n3532), .CLK(clk_in), .RSTB(n7163), .Q(
        \FIFO[32][25] ) );
  DFFARX1 \FIFO_reg[32][24]  ( .D(n3531), .CLK(clk_in), .RSTB(n7163), .Q(
        \FIFO[32][24] ) );
  DFFARX1 \FIFO_reg[32][23]  ( .D(n3530), .CLK(clk_in), .RSTB(n7164), .Q(
        \FIFO[32][23] ) );
  DFFARX1 \FIFO_reg[32][22]  ( .D(n3529), .CLK(clk_in), .RSTB(n7164), .Q(
        \FIFO[32][22] ) );
  DFFARX1 \FIFO_reg[32][21]  ( .D(n3528), .CLK(clk_in), .RSTB(n7164), .Q(
        \FIFO[32][21] ) );
  DFFARX1 \FIFO_reg[32][20]  ( .D(n3527), .CLK(clk_in), .RSTB(n7164), .Q(
        \FIFO[32][20] ) );
  DFFARX1 \FIFO_reg[32][19]  ( .D(n3526), .CLK(clk_in), .RSTB(n7164), .Q(
        \FIFO[32][19] ) );
  DFFARX1 \FIFO_reg[32][18]  ( .D(n3525), .CLK(clk_in), .RSTB(n7164), .Q(
        \FIFO[32][18] ) );
  DFFARX1 \FIFO_reg[32][17]  ( .D(n3524), .CLK(clk_in), .RSTB(n7164), .Q(
        \FIFO[32][17] ) );
  DFFARX1 \FIFO_reg[32][16]  ( .D(n3523), .CLK(clk_in), .RSTB(n7164), .Q(
        \FIFO[32][16] ) );
  DFFARX1 \FIFO_reg[32][15]  ( .D(n3522), .CLK(clk_in), .RSTB(n7164), .Q(
        \FIFO[32][15] ) );
  DFFARX1 \FIFO_reg[32][14]  ( .D(n3521), .CLK(clk_in), .RSTB(n7164), .Q(
        \FIFO[32][14] ) );
  DFFARX1 \FIFO_reg[32][13]  ( .D(n3520), .CLK(clk_in), .RSTB(n7164), .Q(
        \FIFO[32][13] ) );
  DFFARX1 \FIFO_reg[32][12]  ( .D(n3519), .CLK(clk_in), .RSTB(n7164), .Q(
        \FIFO[32][12] ) );
  DFFARX1 \FIFO_reg[32][11]  ( .D(n3518), .CLK(clk_in), .RSTB(n7164), .Q(
        \FIFO[32][11] ) );
  DFFARX1 \FIFO_reg[32][10]  ( .D(n3517), .CLK(clk_in), .RSTB(n7164), .Q(
        \FIFO[32][10] ) );
  DFFARX1 \FIFO_reg[32][9]  ( .D(n3516), .CLK(clk_in), .RSTB(n7164), .Q(
        \FIFO[32][9] ) );
  DFFARX1 \FIFO_reg[32][8]  ( .D(n3515), .CLK(clk_in), .RSTB(n7164), .Q(
        \FIFO[32][8] ) );
  DFFARX1 \FIFO_reg[32][7]  ( .D(n3514), .CLK(clk_in), .RSTB(n7164), .Q(
        \FIFO[32][7] ) );
  DFFARX1 \FIFO_reg[32][6]  ( .D(n3513), .CLK(clk_in), .RSTB(n7164), .Q(
        \FIFO[32][6] ) );
  DFFARX1 \FIFO_reg[32][5]  ( .D(n3512), .CLK(clk_in), .RSTB(n7165), .Q(
        \FIFO[32][5] ) );
  DFFARX1 \FIFO_reg[32][4]  ( .D(n3511), .CLK(clk_in), .RSTB(n7165), .Q(
        \FIFO[32][4] ) );
  DFFARX1 \FIFO_reg[32][3]  ( .D(n3510), .CLK(clk_in), .RSTB(n7165), .Q(
        \FIFO[32][3] ) );
  DFFARX1 \FIFO_reg[32][2]  ( .D(n3509), .CLK(clk_in), .RSTB(n7165), .Q(
        \FIFO[32][2] ) );
  DFFARX1 \FIFO_reg[32][1]  ( .D(n3508), .CLK(clk_in), .RSTB(n7165), .Q(
        \FIFO[32][1] ) );
  DFFARX1 \FIFO_reg[32][0]  ( .D(n3507), .CLK(clk_in), .RSTB(n7165), .Q(
        \FIFO[32][0] ) );
  DFFARX1 \FIFO_reg[33][31]  ( .D(n3506), .CLK(clk_in), .RSTB(n7165), .Q(
        \FIFO[33][31] ) );
  DFFARX1 \FIFO_reg[33][30]  ( .D(n3505), .CLK(clk_in), .RSTB(n7165), .Q(
        \FIFO[33][30] ) );
  DFFARX1 \FIFO_reg[33][29]  ( .D(n3504), .CLK(clk_in), .RSTB(n7165), .Q(
        \FIFO[33][29] ) );
  DFFARX1 \FIFO_reg[33][28]  ( .D(n3503), .CLK(clk_in), .RSTB(n7165), .Q(
        \FIFO[33][28] ) );
  DFFARX1 \FIFO_reg[33][27]  ( .D(n3502), .CLK(clk_in), .RSTB(n7165), .Q(
        \FIFO[33][27] ) );
  DFFARX1 \FIFO_reg[33][26]  ( .D(n3501), .CLK(clk_in), .RSTB(n7165), .Q(
        \FIFO[33][26] ) );
  DFFARX1 \FIFO_reg[33][25]  ( .D(n3500), .CLK(clk_in), .RSTB(n7165), .Q(
        \FIFO[33][25] ) );
  DFFARX1 \FIFO_reg[33][24]  ( .D(n3499), .CLK(clk_in), .RSTB(n7165), .Q(
        \FIFO[33][24] ) );
  DFFARX1 \FIFO_reg[33][23]  ( .D(n3498), .CLK(clk_in), .RSTB(n7165), .Q(
        \FIFO[33][23] ) );
  DFFARX1 \FIFO_reg[33][22]  ( .D(n3497), .CLK(clk_in), .RSTB(n7165), .Q(
        \FIFO[33][22] ) );
  DFFARX1 \FIFO_reg[33][21]  ( .D(n3496), .CLK(clk_in), .RSTB(n7165), .Q(
        \FIFO[33][21] ) );
  DFFARX1 \FIFO_reg[33][20]  ( .D(n3495), .CLK(clk_in), .RSTB(n7165), .Q(
        \FIFO[33][20] ) );
  DFFARX1 \FIFO_reg[33][19]  ( .D(n3494), .CLK(clk_in), .RSTB(n7166), .Q(
        \FIFO[33][19] ) );
  DFFARX1 \FIFO_reg[33][18]  ( .D(n3493), .CLK(clk_in), .RSTB(n7166), .Q(
        \FIFO[33][18] ) );
  DFFARX1 \FIFO_reg[33][17]  ( .D(n3492), .CLK(clk_in), .RSTB(n7166), .Q(
        \FIFO[33][17] ) );
  DFFARX1 \FIFO_reg[33][16]  ( .D(n3491), .CLK(clk_in), .RSTB(n7166), .Q(
        \FIFO[33][16] ) );
  DFFARX1 \FIFO_reg[33][15]  ( .D(n3490), .CLK(clk_in), .RSTB(n7166), .Q(
        \FIFO[33][15] ) );
  DFFARX1 \FIFO_reg[33][14]  ( .D(n3489), .CLK(clk_in), .RSTB(n7166), .Q(
        \FIFO[33][14] ) );
  DFFARX1 \FIFO_reg[33][13]  ( .D(n3488), .CLK(clk_in), .RSTB(n7166), .Q(
        \FIFO[33][13] ) );
  DFFARX1 \FIFO_reg[33][12]  ( .D(n3487), .CLK(clk_in), .RSTB(n7166), .Q(
        \FIFO[33][12] ) );
  DFFARX1 \FIFO_reg[33][11]  ( .D(n3486), .CLK(clk_in), .RSTB(n7166), .Q(
        \FIFO[33][11] ) );
  DFFARX1 \FIFO_reg[33][10]  ( .D(n3485), .CLK(clk_in), .RSTB(n7166), .Q(
        \FIFO[33][10] ) );
  DFFARX1 \FIFO_reg[33][9]  ( .D(n3484), .CLK(clk_in), .RSTB(n7166), .Q(
        \FIFO[33][9] ) );
  DFFARX1 \FIFO_reg[33][8]  ( .D(n3483), .CLK(clk_in), .RSTB(n7166), .Q(
        \FIFO[33][8] ) );
  DFFARX1 \FIFO_reg[33][7]  ( .D(n3482), .CLK(clk_in), .RSTB(n7166), .Q(
        \FIFO[33][7] ) );
  DFFARX1 \FIFO_reg[33][6]  ( .D(n3481), .CLK(clk_in), .RSTB(n7166), .Q(
        \FIFO[33][6] ) );
  DFFARX1 \FIFO_reg[33][5]  ( .D(n3480), .CLK(clk_in), .RSTB(n7166), .Q(
        \FIFO[33][5] ) );
  DFFARX1 \FIFO_reg[33][4]  ( .D(n3479), .CLK(clk_in), .RSTB(n7166), .Q(
        \FIFO[33][4] ) );
  DFFARX1 \FIFO_reg[33][3]  ( .D(n3478), .CLK(clk_in), .RSTB(n7166), .Q(
        \FIFO[33][3] ) );
  DFFARX1 \FIFO_reg[33][2]  ( .D(n3477), .CLK(clk_in), .RSTB(n7166), .Q(
        \FIFO[33][2] ) );
  DFFARX1 \FIFO_reg[33][1]  ( .D(n3476), .CLK(clk_in), .RSTB(n7167), .Q(
        \FIFO[33][1] ) );
  DFFARX1 \FIFO_reg[33][0]  ( .D(n3475), .CLK(clk_in), .RSTB(n7167), .Q(
        \FIFO[33][0] ) );
  DFFARX1 \FIFO_reg[34][31]  ( .D(n3474), .CLK(clk_in), .RSTB(n7167), .Q(
        \FIFO[34][31] ) );
  DFFARX1 \FIFO_reg[34][30]  ( .D(n3473), .CLK(clk_in), .RSTB(n7167), .Q(
        \FIFO[34][30] ) );
  DFFARX1 \FIFO_reg[34][29]  ( .D(n3472), .CLK(clk_in), .RSTB(n7167), .Q(
        \FIFO[34][29] ) );
  DFFARX1 \FIFO_reg[34][28]  ( .D(n3471), .CLK(clk_in), .RSTB(n7167), .Q(
        \FIFO[34][28] ) );
  DFFARX1 \FIFO_reg[34][27]  ( .D(n3470), .CLK(clk_in), .RSTB(n7167), .Q(
        \FIFO[34][27] ) );
  DFFARX1 \FIFO_reg[34][26]  ( .D(n3469), .CLK(clk_in), .RSTB(n7167), .Q(
        \FIFO[34][26] ) );
  DFFARX1 \FIFO_reg[34][25]  ( .D(n3468), .CLK(clk_in), .RSTB(n7167), .Q(
        \FIFO[34][25] ) );
  DFFARX1 \FIFO_reg[34][24]  ( .D(n3467), .CLK(clk_in), .RSTB(n7167), .Q(
        \FIFO[34][24] ) );
  DFFARX1 \FIFO_reg[34][23]  ( .D(n3466), .CLK(clk_in), .RSTB(n7167), .Q(
        \FIFO[34][23] ) );
  DFFARX1 \FIFO_reg[34][22]  ( .D(n3465), .CLK(clk_in), .RSTB(n7167), .Q(
        \FIFO[34][22] ) );
  DFFARX1 \FIFO_reg[34][21]  ( .D(n3464), .CLK(clk_in), .RSTB(n7167), .Q(
        \FIFO[34][21] ) );
  DFFARX1 \FIFO_reg[34][20]  ( .D(n3463), .CLK(clk_in), .RSTB(n7167), .Q(
        \FIFO[34][20] ) );
  DFFARX1 \FIFO_reg[34][19]  ( .D(n3462), .CLK(clk_in), .RSTB(n7167), .Q(
        \FIFO[34][19] ) );
  DFFARX1 \FIFO_reg[34][18]  ( .D(n3461), .CLK(clk_in), .RSTB(n7167), .Q(
        \FIFO[34][18] ) );
  DFFARX1 \FIFO_reg[34][17]  ( .D(n3460), .CLK(clk_in), .RSTB(n7167), .Q(
        \FIFO[34][17] ) );
  DFFARX1 \FIFO_reg[34][16]  ( .D(n3459), .CLK(clk_in), .RSTB(n7167), .Q(
        \FIFO[34][16] ) );
  DFFARX1 \FIFO_reg[34][15]  ( .D(n3458), .CLK(clk_in), .RSTB(n7168), .Q(
        \FIFO[34][15] ) );
  DFFARX1 \FIFO_reg[34][14]  ( .D(n3457), .CLK(clk_in), .RSTB(n7168), .Q(
        \FIFO[34][14] ) );
  DFFARX1 \FIFO_reg[34][13]  ( .D(n3456), .CLK(clk_in), .RSTB(n7168), .Q(
        \FIFO[34][13] ) );
  DFFARX1 \FIFO_reg[34][12]  ( .D(n3455), .CLK(clk_in), .RSTB(n7168), .Q(
        \FIFO[34][12] ) );
  DFFARX1 \FIFO_reg[34][11]  ( .D(n3454), .CLK(clk_in), .RSTB(n7168), .Q(
        \FIFO[34][11] ) );
  DFFARX1 \FIFO_reg[34][10]  ( .D(n3453), .CLK(clk_in), .RSTB(n7168), .Q(
        \FIFO[34][10] ) );
  DFFARX1 \FIFO_reg[34][9]  ( .D(n3452), .CLK(clk_in), .RSTB(n7168), .Q(
        \FIFO[34][9] ) );
  DFFARX1 \FIFO_reg[34][8]  ( .D(n3451), .CLK(clk_in), .RSTB(n7168), .Q(
        \FIFO[34][8] ) );
  DFFARX1 \FIFO_reg[34][7]  ( .D(n3450), .CLK(clk_in), .RSTB(n7168), .Q(
        \FIFO[34][7] ) );
  DFFARX1 \FIFO_reg[34][6]  ( .D(n3449), .CLK(clk_in), .RSTB(n7168), .Q(
        \FIFO[34][6] ) );
  DFFARX1 \FIFO_reg[34][5]  ( .D(n3448), .CLK(clk_in), .RSTB(n7168), .Q(
        \FIFO[34][5] ) );
  DFFARX1 \FIFO_reg[34][4]  ( .D(n3447), .CLK(clk_in), .RSTB(n7168), .Q(
        \FIFO[34][4] ) );
  DFFARX1 \FIFO_reg[34][3]  ( .D(n3446), .CLK(clk_in), .RSTB(n7168), .Q(
        \FIFO[34][3] ) );
  DFFARX1 \FIFO_reg[34][2]  ( .D(n3445), .CLK(clk_in), .RSTB(n7168), .Q(
        \FIFO[34][2] ) );
  DFFARX1 \FIFO_reg[34][1]  ( .D(n3444), .CLK(clk_in), .RSTB(n7168), .Q(
        \FIFO[34][1] ) );
  DFFARX1 \FIFO_reg[34][0]  ( .D(n3443), .CLK(clk_in), .RSTB(n7168), .Q(
        \FIFO[34][0] ) );
  DFFARX1 \FIFO_reg[35][31]  ( .D(n3442), .CLK(clk_in), .RSTB(n7168), .Q(
        \FIFO[35][31] ) );
  DFFARX1 \FIFO_reg[35][30]  ( .D(n3441), .CLK(clk_in), .RSTB(n7168), .Q(
        \FIFO[35][30] ) );
  DFFARX1 \FIFO_reg[35][29]  ( .D(n3440), .CLK(clk_in), .RSTB(n7169), .Q(
        \FIFO[35][29] ) );
  DFFARX1 \FIFO_reg[35][28]  ( .D(n3439), .CLK(clk_in), .RSTB(n7169), .Q(
        \FIFO[35][28] ) );
  DFFARX1 \FIFO_reg[35][27]  ( .D(n3438), .CLK(clk_in), .RSTB(n7169), .Q(
        \FIFO[35][27] ) );
  DFFARX1 \FIFO_reg[35][26]  ( .D(n3437), .CLK(clk_in), .RSTB(n7169), .Q(
        \FIFO[35][26] ) );
  DFFARX1 \FIFO_reg[35][25]  ( .D(n3436), .CLK(clk_in), .RSTB(n7169), .Q(
        \FIFO[35][25] ) );
  DFFARX1 \FIFO_reg[35][24]  ( .D(n3435), .CLK(clk_in), .RSTB(n7169), .Q(
        \FIFO[35][24] ) );
  DFFARX1 \FIFO_reg[35][23]  ( .D(n3434), .CLK(clk_in), .RSTB(n7169), .Q(
        \FIFO[35][23] ) );
  DFFARX1 \FIFO_reg[35][22]  ( .D(n3433), .CLK(clk_in), .RSTB(n7169), .Q(
        \FIFO[35][22] ) );
  DFFARX1 \FIFO_reg[35][21]  ( .D(n3432), .CLK(clk_in), .RSTB(n7169), .Q(
        \FIFO[35][21] ) );
  DFFARX1 \FIFO_reg[35][20]  ( .D(n3431), .CLK(clk_in), .RSTB(n7169), .Q(
        \FIFO[35][20] ) );
  DFFARX1 \FIFO_reg[35][19]  ( .D(n3430), .CLK(clk_in), .RSTB(n7169), .Q(
        \FIFO[35][19] ) );
  DFFARX1 \FIFO_reg[35][18]  ( .D(n3429), .CLK(clk_in), .RSTB(n7169), .Q(
        \FIFO[35][18] ) );
  DFFARX1 \FIFO_reg[35][17]  ( .D(n3428), .CLK(clk_in), .RSTB(n7169), .Q(
        \FIFO[35][17] ) );
  DFFARX1 \FIFO_reg[35][16]  ( .D(n3427), .CLK(clk_in), .RSTB(n7169), .Q(
        \FIFO[35][16] ) );
  DFFARX1 \FIFO_reg[35][15]  ( .D(n3426), .CLK(clk_in), .RSTB(n7169), .Q(
        \FIFO[35][15] ) );
  DFFARX1 \FIFO_reg[35][14]  ( .D(n3425), .CLK(clk_in), .RSTB(n7169), .Q(
        \FIFO[35][14] ) );
  DFFARX1 \FIFO_reg[35][13]  ( .D(n3424), .CLK(clk_in), .RSTB(n7169), .Q(
        \FIFO[35][13] ) );
  DFFARX1 \FIFO_reg[35][12]  ( .D(n3423), .CLK(clk_in), .RSTB(n7169), .Q(
        \FIFO[35][12] ) );
  DFFARX1 \FIFO_reg[35][11]  ( .D(n3422), .CLK(clk_in), .RSTB(n7170), .Q(
        \FIFO[35][11] ) );
  DFFARX1 \FIFO_reg[35][10]  ( .D(n3421), .CLK(clk_in), .RSTB(n7170), .Q(
        \FIFO[35][10] ) );
  DFFARX1 \FIFO_reg[35][9]  ( .D(n3420), .CLK(clk_in), .RSTB(n7170), .Q(
        \FIFO[35][9] ) );
  DFFARX1 \FIFO_reg[35][8]  ( .D(n3419), .CLK(clk_in), .RSTB(n7170), .Q(
        \FIFO[35][8] ) );
  DFFARX1 \FIFO_reg[35][7]  ( .D(n3418), .CLK(clk_in), .RSTB(n7170), .Q(
        \FIFO[35][7] ) );
  DFFARX1 \FIFO_reg[35][6]  ( .D(n3417), .CLK(clk_in), .RSTB(n7170), .Q(
        \FIFO[35][6] ) );
  DFFARX1 \FIFO_reg[35][5]  ( .D(n3416), .CLK(clk_in), .RSTB(n7170), .Q(
        \FIFO[35][5] ) );
  DFFARX1 \FIFO_reg[35][4]  ( .D(n3415), .CLK(clk_in), .RSTB(n7170), .Q(
        \FIFO[35][4] ) );
  DFFARX1 \FIFO_reg[35][3]  ( .D(n3414), .CLK(clk_in), .RSTB(n7170), .Q(
        \FIFO[35][3] ) );
  DFFARX1 \FIFO_reg[35][2]  ( .D(n3413), .CLK(clk_in), .RSTB(n7170), .Q(
        \FIFO[35][2] ) );
  DFFARX1 \FIFO_reg[35][1]  ( .D(n3412), .CLK(clk_in), .RSTB(n7170), .Q(
        \FIFO[35][1] ) );
  DFFARX1 \FIFO_reg[35][0]  ( .D(n3411), .CLK(clk_in), .RSTB(n7170), .Q(
        \FIFO[35][0] ) );
  DFFARX1 \FIFO_reg[36][31]  ( .D(n3410), .CLK(clk_in), .RSTB(n7170), .Q(
        \FIFO[36][31] ) );
  DFFARX1 \FIFO_reg[36][30]  ( .D(n3409), .CLK(clk_in), .RSTB(n7170), .Q(
        \FIFO[36][30] ) );
  DFFARX1 \FIFO_reg[36][29]  ( .D(n3408), .CLK(clk_in), .RSTB(n7170), .Q(
        \FIFO[36][29] ) );
  DFFARX1 \FIFO_reg[36][28]  ( .D(n3407), .CLK(clk_in), .RSTB(n7170), .Q(
        \FIFO[36][28] ) );
  DFFARX1 \FIFO_reg[36][27]  ( .D(n3406), .CLK(clk_in), .RSTB(n7170), .Q(
        \FIFO[36][27] ) );
  DFFARX1 \FIFO_reg[36][26]  ( .D(n3405), .CLK(clk_in), .RSTB(n7170), .Q(
        \FIFO[36][26] ) );
  DFFARX1 \FIFO_reg[36][25]  ( .D(n3404), .CLK(clk_in), .RSTB(n7171), .Q(
        \FIFO[36][25] ) );
  DFFARX1 \FIFO_reg[36][24]  ( .D(n3403), .CLK(clk_in), .RSTB(n7171), .Q(
        \FIFO[36][24] ) );
  DFFARX1 \FIFO_reg[36][23]  ( .D(n3402), .CLK(clk_in), .RSTB(n7171), .Q(
        \FIFO[36][23] ) );
  DFFARX1 \FIFO_reg[36][22]  ( .D(n3401), .CLK(clk_in), .RSTB(n7171), .Q(
        \FIFO[36][22] ) );
  DFFARX1 \FIFO_reg[36][21]  ( .D(n3400), .CLK(clk_in), .RSTB(n7171), .Q(
        \FIFO[36][21] ) );
  DFFARX1 \FIFO_reg[36][20]  ( .D(n3399), .CLK(clk_in), .RSTB(n7171), .Q(
        \FIFO[36][20] ) );
  DFFARX1 \FIFO_reg[36][19]  ( .D(n3398), .CLK(clk_in), .RSTB(n7171), .Q(
        \FIFO[36][19] ) );
  DFFARX1 \FIFO_reg[36][18]  ( .D(n3397), .CLK(clk_in), .RSTB(n7171), .Q(
        \FIFO[36][18] ) );
  DFFARX1 \FIFO_reg[36][17]  ( .D(n3396), .CLK(clk_in), .RSTB(n7171), .Q(
        \FIFO[36][17] ) );
  DFFARX1 \FIFO_reg[36][16]  ( .D(n3395), .CLK(clk_in), .RSTB(n7171), .Q(
        \FIFO[36][16] ) );
  DFFARX1 \FIFO_reg[36][15]  ( .D(n3394), .CLK(clk_in), .RSTB(n7171), .Q(
        \FIFO[36][15] ) );
  DFFARX1 \FIFO_reg[36][14]  ( .D(n3393), .CLK(clk_in), .RSTB(n7171), .Q(
        \FIFO[36][14] ) );
  DFFARX1 \FIFO_reg[36][13]  ( .D(n3392), .CLK(clk_in), .RSTB(n7171), .Q(
        \FIFO[36][13] ) );
  DFFARX1 \FIFO_reg[36][12]  ( .D(n3391), .CLK(clk_in), .RSTB(n7171), .Q(
        \FIFO[36][12] ) );
  DFFARX1 \FIFO_reg[36][11]  ( .D(n3390), .CLK(clk_in), .RSTB(n7171), .Q(
        \FIFO[36][11] ) );
  DFFARX1 \FIFO_reg[36][10]  ( .D(n3389), .CLK(clk_in), .RSTB(n7171), .Q(
        \FIFO[36][10] ) );
  DFFARX1 \FIFO_reg[36][9]  ( .D(n3388), .CLK(clk_in), .RSTB(n7171), .Q(
        \FIFO[36][9] ) );
  DFFARX1 \FIFO_reg[36][8]  ( .D(n3387), .CLK(clk_in), .RSTB(n7171), .Q(
        \FIFO[36][8] ) );
  DFFARX1 \FIFO_reg[36][7]  ( .D(n3386), .CLK(clk_in), .RSTB(n7172), .Q(
        \FIFO[36][7] ) );
  DFFARX1 \FIFO_reg[36][6]  ( .D(n3385), .CLK(clk_in), .RSTB(n7172), .Q(
        \FIFO[36][6] ) );
  DFFARX1 \FIFO_reg[36][5]  ( .D(n3384), .CLK(clk_in), .RSTB(n7172), .Q(
        \FIFO[36][5] ) );
  DFFARX1 \FIFO_reg[36][4]  ( .D(n3383), .CLK(clk_in), .RSTB(n7172), .Q(
        \FIFO[36][4] ) );
  DFFARX1 \FIFO_reg[36][3]  ( .D(n3382), .CLK(clk_in), .RSTB(n7172), .Q(
        \FIFO[36][3] ) );
  DFFARX1 \FIFO_reg[36][2]  ( .D(n3381), .CLK(clk_in), .RSTB(n7172), .Q(
        \FIFO[36][2] ) );
  DFFARX1 \FIFO_reg[36][1]  ( .D(n3380), .CLK(clk_in), .RSTB(n7172), .Q(
        \FIFO[36][1] ) );
  DFFARX1 \FIFO_reg[36][0]  ( .D(n3379), .CLK(clk_in), .RSTB(n7172), .Q(
        \FIFO[36][0] ) );
  DFFARX1 \FIFO_reg[37][31]  ( .D(n3378), .CLK(clk_in), .RSTB(n7172), .Q(
        \FIFO[37][31] ) );
  DFFARX1 \FIFO_reg[37][30]  ( .D(n3377), .CLK(clk_in), .RSTB(n7172), .Q(
        \FIFO[37][30] ) );
  DFFARX1 \FIFO_reg[37][29]  ( .D(n3376), .CLK(clk_in), .RSTB(n7172), .Q(
        \FIFO[37][29] ) );
  DFFARX1 \FIFO_reg[37][28]  ( .D(n3375), .CLK(clk_in), .RSTB(n7172), .Q(
        \FIFO[37][28] ) );
  DFFARX1 \FIFO_reg[37][27]  ( .D(n3374), .CLK(clk_in), .RSTB(n7172), .Q(
        \FIFO[37][27] ) );
  DFFARX1 \FIFO_reg[37][26]  ( .D(n3373), .CLK(clk_in), .RSTB(n7172), .Q(
        \FIFO[37][26] ) );
  DFFARX1 \FIFO_reg[37][25]  ( .D(n3372), .CLK(clk_in), .RSTB(n7172), .Q(
        \FIFO[37][25] ) );
  DFFARX1 \FIFO_reg[37][24]  ( .D(n3371), .CLK(clk_in), .RSTB(n7172), .Q(
        \FIFO[37][24] ) );
  DFFARX1 \FIFO_reg[37][23]  ( .D(n3370), .CLK(clk_in), .RSTB(n7172), .Q(
        \FIFO[37][23] ) );
  DFFARX1 \FIFO_reg[37][22]  ( .D(n3369), .CLK(clk_in), .RSTB(n7172), .Q(
        \FIFO[37][22] ) );
  DFFARX1 \FIFO_reg[37][21]  ( .D(n3368), .CLK(clk_in), .RSTB(n7173), .Q(
        \FIFO[37][21] ) );
  DFFARX1 \FIFO_reg[37][20]  ( .D(n3367), .CLK(clk_in), .RSTB(n7173), .Q(
        \FIFO[37][20] ) );
  DFFARX1 \FIFO_reg[37][19]  ( .D(n3366), .CLK(clk_in), .RSTB(n7173), .Q(
        \FIFO[37][19] ) );
  DFFARX1 \FIFO_reg[37][18]  ( .D(n3365), .CLK(clk_in), .RSTB(n7173), .Q(
        \FIFO[37][18] ) );
  DFFARX1 \FIFO_reg[37][17]  ( .D(n3364), .CLK(clk_in), .RSTB(n7173), .Q(
        \FIFO[37][17] ) );
  DFFARX1 \FIFO_reg[37][16]  ( .D(n3363), .CLK(clk_in), .RSTB(n7173), .Q(
        \FIFO[37][16] ) );
  DFFARX1 \FIFO_reg[37][15]  ( .D(n3362), .CLK(clk_in), .RSTB(n7173), .Q(
        \FIFO[37][15] ) );
  DFFARX1 \FIFO_reg[37][14]  ( .D(n3361), .CLK(clk_in), .RSTB(n7173), .Q(
        \FIFO[37][14] ) );
  DFFARX1 \FIFO_reg[37][13]  ( .D(n3360), .CLK(clk_in), .RSTB(n7173), .Q(
        \FIFO[37][13] ) );
  DFFARX1 \FIFO_reg[37][12]  ( .D(n3359), .CLK(clk_in), .RSTB(n7173), .Q(
        \FIFO[37][12] ) );
  DFFARX1 \FIFO_reg[37][11]  ( .D(n3358), .CLK(clk_in), .RSTB(n7173), .Q(
        \FIFO[37][11] ) );
  DFFARX1 \FIFO_reg[37][10]  ( .D(n3357), .CLK(clk_in), .RSTB(n7173), .Q(
        \FIFO[37][10] ) );
  DFFARX1 \FIFO_reg[37][9]  ( .D(n3356), .CLK(clk_in), .RSTB(n7173), .Q(
        \FIFO[37][9] ) );
  DFFARX1 \FIFO_reg[37][8]  ( .D(n3355), .CLK(clk_in), .RSTB(n7173), .Q(
        \FIFO[37][8] ) );
  DFFARX1 \FIFO_reg[37][7]  ( .D(n3354), .CLK(clk_in), .RSTB(n7173), .Q(
        \FIFO[37][7] ) );
  DFFARX1 \FIFO_reg[37][6]  ( .D(n3353), .CLK(clk_in), .RSTB(n7173), .Q(
        \FIFO[37][6] ) );
  DFFARX1 \FIFO_reg[37][5]  ( .D(n3352), .CLK(clk_in), .RSTB(n7173), .Q(
        \FIFO[37][5] ) );
  DFFARX1 \FIFO_reg[37][4]  ( .D(n3351), .CLK(clk_in), .RSTB(n7173), .Q(
        \FIFO[37][4] ) );
  DFFARX1 \FIFO_reg[37][3]  ( .D(n3350), .CLK(clk_in), .RSTB(n7174), .Q(
        \FIFO[37][3] ) );
  DFFARX1 \FIFO_reg[37][2]  ( .D(n3349), .CLK(clk_in), .RSTB(n7174), .Q(
        \FIFO[37][2] ) );
  DFFARX1 \FIFO_reg[37][1]  ( .D(n3348), .CLK(clk_in), .RSTB(n7174), .Q(
        \FIFO[37][1] ) );
  DFFARX1 \FIFO_reg[37][0]  ( .D(n3347), .CLK(clk_in), .RSTB(n7174), .Q(
        \FIFO[37][0] ) );
  DFFARX1 \FIFO_reg[38][31]  ( .D(n3346), .CLK(clk_in), .RSTB(n7174), .Q(
        \FIFO[38][31] ) );
  DFFARX1 \FIFO_reg[38][30]  ( .D(n3345), .CLK(clk_in), .RSTB(n7174), .Q(
        \FIFO[38][30] ) );
  DFFARX1 \FIFO_reg[38][29]  ( .D(n3344), .CLK(clk_in), .RSTB(n7174), .Q(
        \FIFO[38][29] ) );
  DFFARX1 \FIFO_reg[38][28]  ( .D(n3343), .CLK(clk_in), .RSTB(n7174), .Q(
        \FIFO[38][28] ) );
  DFFARX1 \FIFO_reg[38][27]  ( .D(n3342), .CLK(clk_in), .RSTB(n7174), .Q(
        \FIFO[38][27] ) );
  DFFARX1 \FIFO_reg[38][26]  ( .D(n3341), .CLK(clk_in), .RSTB(n7174), .Q(
        \FIFO[38][26] ) );
  DFFARX1 \FIFO_reg[38][25]  ( .D(n3340), .CLK(clk_in), .RSTB(n7174), .Q(
        \FIFO[38][25] ) );
  DFFARX1 \FIFO_reg[38][24]  ( .D(n3339), .CLK(clk_in), .RSTB(n7174), .Q(
        \FIFO[38][24] ) );
  DFFARX1 \FIFO_reg[38][23]  ( .D(n3338), .CLK(clk_in), .RSTB(n7174), .Q(
        \FIFO[38][23] ) );
  DFFARX1 \FIFO_reg[38][22]  ( .D(n3337), .CLK(clk_in), .RSTB(n7174), .Q(
        \FIFO[38][22] ) );
  DFFARX1 \FIFO_reg[38][21]  ( .D(n3336), .CLK(clk_in), .RSTB(n7174), .Q(
        \FIFO[38][21] ) );
  DFFARX1 \FIFO_reg[38][20]  ( .D(n3335), .CLK(clk_in), .RSTB(n7174), .Q(
        \FIFO[38][20] ) );
  DFFARX1 \FIFO_reg[38][19]  ( .D(n3334), .CLK(clk_in), .RSTB(n7174), .Q(
        \FIFO[38][19] ) );
  DFFARX1 \FIFO_reg[38][18]  ( .D(n3333), .CLK(clk_in), .RSTB(n7174), .Q(
        \FIFO[38][18] ) );
  DFFARX1 \FIFO_reg[38][17]  ( .D(n3332), .CLK(clk_in), .RSTB(n7175), .Q(
        \FIFO[38][17] ) );
  DFFARX1 \FIFO_reg[38][16]  ( .D(n3331), .CLK(clk_in), .RSTB(n7175), .Q(
        \FIFO[38][16] ) );
  DFFARX1 \FIFO_reg[38][15]  ( .D(n3330), .CLK(clk_in), .RSTB(n7175), .Q(
        \FIFO[38][15] ) );
  DFFARX1 \FIFO_reg[38][14]  ( .D(n3329), .CLK(clk_in), .RSTB(n7175), .Q(
        \FIFO[38][14] ) );
  DFFARX1 \FIFO_reg[38][13]  ( .D(n3328), .CLK(clk_in), .RSTB(n7175), .Q(
        \FIFO[38][13] ) );
  DFFARX1 \FIFO_reg[38][12]  ( .D(n3327), .CLK(clk_in), .RSTB(n7175), .Q(
        \FIFO[38][12] ) );
  DFFARX1 \FIFO_reg[38][11]  ( .D(n3326), .CLK(clk_in), .RSTB(n7175), .Q(
        \FIFO[38][11] ) );
  DFFARX1 \FIFO_reg[38][10]  ( .D(n3325), .CLK(clk_in), .RSTB(n7175), .Q(
        \FIFO[38][10] ) );
  DFFARX1 \FIFO_reg[38][9]  ( .D(n3324), .CLK(clk_in), .RSTB(n7175), .Q(
        \FIFO[38][9] ) );
  DFFARX1 \FIFO_reg[38][8]  ( .D(n3323), .CLK(clk_in), .RSTB(n7175), .Q(
        \FIFO[38][8] ) );
  DFFARX1 \FIFO_reg[38][7]  ( .D(n3322), .CLK(clk_in), .RSTB(n7175), .Q(
        \FIFO[38][7] ) );
  DFFARX1 \FIFO_reg[38][6]  ( .D(n3321), .CLK(clk_in), .RSTB(n7175), .Q(
        \FIFO[38][6] ) );
  DFFARX1 \FIFO_reg[38][5]  ( .D(n3320), .CLK(clk_in), .RSTB(n7175), .Q(
        \FIFO[38][5] ) );
  DFFARX1 \FIFO_reg[38][4]  ( .D(n3319), .CLK(clk_in), .RSTB(n7175), .Q(
        \FIFO[38][4] ) );
  DFFARX1 \FIFO_reg[38][3]  ( .D(n3318), .CLK(clk_in), .RSTB(n7175), .Q(
        \FIFO[38][3] ) );
  DFFARX1 \FIFO_reg[38][2]  ( .D(n3317), .CLK(clk_in), .RSTB(n7175), .Q(
        \FIFO[38][2] ) );
  DFFARX1 \FIFO_reg[38][1]  ( .D(n3316), .CLK(clk_in), .RSTB(n7175), .Q(
        \FIFO[38][1] ) );
  DFFARX1 \FIFO_reg[38][0]  ( .D(n3315), .CLK(clk_in), .RSTB(n7175), .Q(
        \FIFO[38][0] ) );
  DFFARX1 \FIFO_reg[39][31]  ( .D(n3314), .CLK(clk_in), .RSTB(n7176), .Q(
        \FIFO[39][31] ) );
  DFFARX1 \FIFO_reg[39][30]  ( .D(n3313), .CLK(clk_in), .RSTB(n7176), .Q(
        \FIFO[39][30] ) );
  DFFARX1 \FIFO_reg[39][29]  ( .D(n3312), .CLK(clk_in), .RSTB(n7176), .Q(
        \FIFO[39][29] ) );
  DFFARX1 \FIFO_reg[39][28]  ( .D(n3311), .CLK(clk_in), .RSTB(n7176), .Q(
        \FIFO[39][28] ) );
  DFFARX1 \FIFO_reg[39][27]  ( .D(n3310), .CLK(clk_in), .RSTB(n7176), .Q(
        \FIFO[39][27] ) );
  DFFARX1 \FIFO_reg[39][26]  ( .D(n3309), .CLK(clk_in), .RSTB(n7176), .Q(
        \FIFO[39][26] ) );
  DFFARX1 \FIFO_reg[39][25]  ( .D(n3308), .CLK(clk_in), .RSTB(n7176), .Q(
        \FIFO[39][25] ) );
  DFFARX1 \FIFO_reg[39][24]  ( .D(n3307), .CLK(clk_in), .RSTB(n7176), .Q(
        \FIFO[39][24] ) );
  DFFARX1 \FIFO_reg[39][23]  ( .D(n3306), .CLK(clk_in), .RSTB(n7176), .Q(
        \FIFO[39][23] ) );
  DFFARX1 \FIFO_reg[39][22]  ( .D(n3305), .CLK(clk_in), .RSTB(n7176), .Q(
        \FIFO[39][22] ) );
  DFFARX1 \FIFO_reg[39][21]  ( .D(n3304), .CLK(clk_in), .RSTB(n7176), .Q(
        \FIFO[39][21] ) );
  DFFARX1 \FIFO_reg[39][20]  ( .D(n3303), .CLK(clk_in), .RSTB(n7176), .Q(
        \FIFO[39][20] ) );
  DFFARX1 \FIFO_reg[39][19]  ( .D(n3302), .CLK(clk_in), .RSTB(n7176), .Q(
        \FIFO[39][19] ) );
  DFFARX1 \FIFO_reg[39][18]  ( .D(n3301), .CLK(clk_in), .RSTB(n7176), .Q(
        \FIFO[39][18] ) );
  DFFARX1 \FIFO_reg[39][17]  ( .D(n3300), .CLK(clk_in), .RSTB(n7176), .Q(
        \FIFO[39][17] ) );
  DFFARX1 \FIFO_reg[39][16]  ( .D(n3299), .CLK(clk_in), .RSTB(n7176), .Q(
        \FIFO[39][16] ) );
  DFFARX1 \FIFO_reg[39][15]  ( .D(n3298), .CLK(clk_in), .RSTB(n7176), .Q(
        \FIFO[39][15] ) );
  DFFARX1 \FIFO_reg[39][14]  ( .D(n3297), .CLK(clk_in), .RSTB(n7176), .Q(
        \FIFO[39][14] ) );
  DFFARX1 \FIFO_reg[39][13]  ( .D(n3296), .CLK(clk_in), .RSTB(n7177), .Q(
        \FIFO[39][13] ) );
  DFFARX1 \FIFO_reg[39][12]  ( .D(n3295), .CLK(clk_in), .RSTB(n7177), .Q(
        \FIFO[39][12] ) );
  DFFARX1 \FIFO_reg[39][11]  ( .D(n3294), .CLK(clk_in), .RSTB(n7177), .Q(
        \FIFO[39][11] ) );
  DFFARX1 \FIFO_reg[39][10]  ( .D(n3293), .CLK(clk_in), .RSTB(n7177), .Q(
        \FIFO[39][10] ) );
  DFFARX1 \FIFO_reg[39][9]  ( .D(n3292), .CLK(clk_in), .RSTB(n7177), .Q(
        \FIFO[39][9] ) );
  DFFARX1 \FIFO_reg[39][8]  ( .D(n3291), .CLK(clk_in), .RSTB(n7177), .Q(
        \FIFO[39][8] ) );
  DFFARX1 \FIFO_reg[39][7]  ( .D(n3290), .CLK(clk_in), .RSTB(n7177), .Q(
        \FIFO[39][7] ) );
  DFFARX1 \FIFO_reg[39][6]  ( .D(n3289), .CLK(clk_in), .RSTB(n7177), .Q(
        \FIFO[39][6] ) );
  DFFARX1 \FIFO_reg[39][5]  ( .D(n3288), .CLK(clk_in), .RSTB(n7177), .Q(
        \FIFO[39][5] ) );
  DFFARX1 \FIFO_reg[39][4]  ( .D(n3287), .CLK(clk_in), .RSTB(n7177), .Q(
        \FIFO[39][4] ) );
  DFFARX1 \FIFO_reg[39][3]  ( .D(n3286), .CLK(clk_in), .RSTB(n7177), .Q(
        \FIFO[39][3] ) );
  DFFARX1 \FIFO_reg[39][2]  ( .D(n3285), .CLK(clk_in), .RSTB(n7177), .Q(
        \FIFO[39][2] ) );
  DFFARX1 \FIFO_reg[39][1]  ( .D(n3284), .CLK(clk_in), .RSTB(n7177), .Q(
        \FIFO[39][1] ) );
  DFFARX1 \FIFO_reg[39][0]  ( .D(n3283), .CLK(clk_in), .RSTB(n7177), .Q(
        \FIFO[39][0] ) );
  DFFARX1 \FIFO_reg[40][31]  ( .D(n3282), .CLK(clk_in), .RSTB(n7177), .Q(
        \FIFO[40][31] ) );
  DFFARX1 \FIFO_reg[40][30]  ( .D(n3281), .CLK(clk_in), .RSTB(n7177), .Q(
        \FIFO[40][30] ) );
  DFFARX1 \FIFO_reg[40][29]  ( .D(n3280), .CLK(clk_in), .RSTB(n7177), .Q(
        \FIFO[40][29] ) );
  DFFARX1 \FIFO_reg[40][28]  ( .D(n3279), .CLK(clk_in), .RSTB(n7177), .Q(
        \FIFO[40][28] ) );
  DFFARX1 \FIFO_reg[40][27]  ( .D(n3278), .CLK(clk_in), .RSTB(n7178), .Q(
        \FIFO[40][27] ) );
  DFFARX1 \FIFO_reg[40][26]  ( .D(n3277), .CLK(clk_in), .RSTB(n7178), .Q(
        \FIFO[40][26] ) );
  DFFARX1 \FIFO_reg[40][25]  ( .D(n3276), .CLK(clk_in), .RSTB(n7178), .Q(
        \FIFO[40][25] ) );
  DFFARX1 \FIFO_reg[40][24]  ( .D(n3275), .CLK(clk_in), .RSTB(n7178), .Q(
        \FIFO[40][24] ) );
  DFFARX1 \FIFO_reg[40][23]  ( .D(n3274), .CLK(clk_in), .RSTB(n7178), .Q(
        \FIFO[40][23] ) );
  DFFARX1 \FIFO_reg[40][22]  ( .D(n3273), .CLK(clk_in), .RSTB(n7178), .Q(
        \FIFO[40][22] ) );
  DFFARX1 \FIFO_reg[40][21]  ( .D(n3272), .CLK(clk_in), .RSTB(n7178), .Q(
        \FIFO[40][21] ) );
  DFFARX1 \FIFO_reg[40][20]  ( .D(n3271), .CLK(clk_in), .RSTB(n7178), .Q(
        \FIFO[40][20] ) );
  DFFARX1 \FIFO_reg[40][19]  ( .D(n3270), .CLK(clk_in), .RSTB(n7178), .Q(
        \FIFO[40][19] ) );
  DFFARX1 \FIFO_reg[40][18]  ( .D(n3269), .CLK(clk_in), .RSTB(n7178), .Q(
        \FIFO[40][18] ) );
  DFFARX1 \FIFO_reg[40][17]  ( .D(n3268), .CLK(clk_in), .RSTB(n7178), .Q(
        \FIFO[40][17] ) );
  DFFARX1 \FIFO_reg[40][16]  ( .D(n3267), .CLK(clk_in), .RSTB(n7178), .Q(
        \FIFO[40][16] ) );
  DFFARX1 \FIFO_reg[40][15]  ( .D(n3266), .CLK(clk_in), .RSTB(n7178), .Q(
        \FIFO[40][15] ) );
  DFFARX1 \FIFO_reg[40][14]  ( .D(n3265), .CLK(clk_in), .RSTB(n7178), .Q(
        \FIFO[40][14] ) );
  DFFARX1 \FIFO_reg[40][13]  ( .D(n3264), .CLK(clk_in), .RSTB(n7178), .Q(
        \FIFO[40][13] ) );
  DFFARX1 \FIFO_reg[40][12]  ( .D(n3263), .CLK(clk_in), .RSTB(n7178), .Q(
        \FIFO[40][12] ) );
  DFFARX1 \FIFO_reg[40][11]  ( .D(n3262), .CLK(clk_in), .RSTB(n7178), .Q(
        \FIFO[40][11] ) );
  DFFARX1 \FIFO_reg[40][10]  ( .D(n3261), .CLK(clk_in), .RSTB(n7178), .Q(
        \FIFO[40][10] ) );
  DFFARX1 \FIFO_reg[40][9]  ( .D(n3260), .CLK(clk_in), .RSTB(n7179), .Q(
        \FIFO[40][9] ) );
  DFFARX1 \FIFO_reg[40][8]  ( .D(n3259), .CLK(clk_in), .RSTB(n7179), .Q(
        \FIFO[40][8] ) );
  DFFARX1 \FIFO_reg[40][7]  ( .D(n3258), .CLK(clk_in), .RSTB(n7179), .Q(
        \FIFO[40][7] ) );
  DFFARX1 \FIFO_reg[40][6]  ( .D(n3257), .CLK(clk_in), .RSTB(n7179), .Q(
        \FIFO[40][6] ) );
  DFFARX1 \FIFO_reg[40][5]  ( .D(n3256), .CLK(clk_in), .RSTB(n7179), .Q(
        \FIFO[40][5] ) );
  DFFARX1 \FIFO_reg[40][4]  ( .D(n3255), .CLK(clk_in), .RSTB(n7179), .Q(
        \FIFO[40][4] ) );
  DFFARX1 \FIFO_reg[40][3]  ( .D(n3254), .CLK(clk_in), .RSTB(n7179), .Q(
        \FIFO[40][3] ) );
  DFFARX1 \FIFO_reg[40][2]  ( .D(n3253), .CLK(clk_in), .RSTB(n7179), .Q(
        \FIFO[40][2] ) );
  DFFARX1 \FIFO_reg[40][1]  ( .D(n3252), .CLK(clk_in), .RSTB(n7179), .Q(
        \FIFO[40][1] ) );
  DFFARX1 \FIFO_reg[40][0]  ( .D(n3251), .CLK(clk_in), .RSTB(n7179), .Q(
        \FIFO[40][0] ) );
  DFFARX1 \FIFO_reg[41][31]  ( .D(n3250), .CLK(clk_in), .RSTB(n7179), .Q(
        \FIFO[41][31] ) );
  DFFARX1 \FIFO_reg[41][30]  ( .D(n3249), .CLK(clk_in), .RSTB(n7179), .Q(
        \FIFO[41][30] ) );
  DFFARX1 \FIFO_reg[41][29]  ( .D(n3248), .CLK(clk_in), .RSTB(n7179), .Q(
        \FIFO[41][29] ) );
  DFFARX1 \FIFO_reg[41][28]  ( .D(n3247), .CLK(clk_in), .RSTB(n7179), .Q(
        \FIFO[41][28] ) );
  DFFARX1 \FIFO_reg[41][27]  ( .D(n3246), .CLK(clk_in), .RSTB(n7179), .Q(
        \FIFO[41][27] ) );
  DFFARX1 \FIFO_reg[41][26]  ( .D(n3245), .CLK(clk_in), .RSTB(n7179), .Q(
        \FIFO[41][26] ) );
  DFFARX1 \FIFO_reg[41][25]  ( .D(n3244), .CLK(clk_in), .RSTB(n7179), .Q(
        \FIFO[41][25] ) );
  DFFARX1 \FIFO_reg[41][24]  ( .D(n3243), .CLK(clk_in), .RSTB(n7179), .Q(
        \FIFO[41][24] ) );
  DFFARX1 \FIFO_reg[41][23]  ( .D(n3242), .CLK(clk_in), .RSTB(n7180), .Q(
        \FIFO[41][23] ) );
  DFFARX1 \FIFO_reg[41][22]  ( .D(n3241), .CLK(clk_in), .RSTB(n7180), .Q(
        \FIFO[41][22] ) );
  DFFARX1 \FIFO_reg[41][21]  ( .D(n3240), .CLK(clk_in), .RSTB(n7180), .Q(
        \FIFO[41][21] ) );
  DFFARX1 \FIFO_reg[41][20]  ( .D(n3239), .CLK(clk_in), .RSTB(n7180), .Q(
        \FIFO[41][20] ) );
  DFFARX1 \FIFO_reg[41][19]  ( .D(n3238), .CLK(clk_in), .RSTB(n7180), .Q(
        \FIFO[41][19] ) );
  DFFARX1 \FIFO_reg[41][18]  ( .D(n3237), .CLK(clk_in), .RSTB(n7180), .Q(
        \FIFO[41][18] ) );
  DFFARX1 \FIFO_reg[41][17]  ( .D(n3236), .CLK(clk_in), .RSTB(n7180), .Q(
        \FIFO[41][17] ) );
  DFFARX1 \FIFO_reg[41][16]  ( .D(n3235), .CLK(clk_in), .RSTB(n7180), .Q(
        \FIFO[41][16] ) );
  DFFARX1 \FIFO_reg[41][15]  ( .D(n3234), .CLK(clk_in), .RSTB(n7180), .Q(
        \FIFO[41][15] ) );
  DFFARX1 \FIFO_reg[41][14]  ( .D(n3233), .CLK(clk_in), .RSTB(n7180), .Q(
        \FIFO[41][14] ) );
  DFFARX1 \FIFO_reg[41][13]  ( .D(n3232), .CLK(clk_in), .RSTB(n7180), .Q(
        \FIFO[41][13] ) );
  DFFARX1 \FIFO_reg[41][12]  ( .D(n3231), .CLK(clk_in), .RSTB(n7180), .Q(
        \FIFO[41][12] ) );
  DFFARX1 \FIFO_reg[41][11]  ( .D(n3230), .CLK(clk_in), .RSTB(n7180), .Q(
        \FIFO[41][11] ) );
  DFFARX1 \FIFO_reg[41][10]  ( .D(n3229), .CLK(clk_in), .RSTB(n7180), .Q(
        \FIFO[41][10] ) );
  DFFARX1 \FIFO_reg[41][9]  ( .D(n3228), .CLK(clk_in), .RSTB(n7180), .Q(
        \FIFO[41][9] ) );
  DFFARX1 \FIFO_reg[41][8]  ( .D(n3227), .CLK(clk_in), .RSTB(n7180), .Q(
        \FIFO[41][8] ) );
  DFFARX1 \FIFO_reg[41][7]  ( .D(n3226), .CLK(clk_in), .RSTB(n7180), .Q(
        \FIFO[41][7] ) );
  DFFARX1 \FIFO_reg[41][6]  ( .D(n3225), .CLK(clk_in), .RSTB(n7180), .Q(
        \FIFO[41][6] ) );
  DFFARX1 \FIFO_reg[41][5]  ( .D(n3224), .CLK(clk_in), .RSTB(n7181), .Q(
        \FIFO[41][5] ) );
  DFFARX1 \FIFO_reg[41][4]  ( .D(n3223), .CLK(clk_in), .RSTB(n7181), .Q(
        \FIFO[41][4] ) );
  DFFARX1 \FIFO_reg[41][3]  ( .D(n3222), .CLK(clk_in), .RSTB(n7181), .Q(
        \FIFO[41][3] ) );
  DFFARX1 \FIFO_reg[41][2]  ( .D(n3221), .CLK(clk_in), .RSTB(n7181), .Q(
        \FIFO[41][2] ) );
  DFFARX1 \FIFO_reg[41][1]  ( .D(n3220), .CLK(clk_in), .RSTB(n7181), .Q(
        \FIFO[41][1] ) );
  DFFARX1 \FIFO_reg[41][0]  ( .D(n3219), .CLK(clk_in), .RSTB(n7181), .Q(
        \FIFO[41][0] ) );
  DFFARX1 \FIFO_reg[42][31]  ( .D(n3218), .CLK(clk_in), .RSTB(n7181), .Q(
        \FIFO[42][31] ) );
  DFFARX1 \FIFO_reg[42][30]  ( .D(n3217), .CLK(clk_in), .RSTB(n7181), .Q(
        \FIFO[42][30] ) );
  DFFARX1 \FIFO_reg[42][29]  ( .D(n3216), .CLK(clk_in), .RSTB(n7181), .Q(
        \FIFO[42][29] ) );
  DFFARX1 \FIFO_reg[42][28]  ( .D(n3215), .CLK(clk_in), .RSTB(n7181), .Q(
        \FIFO[42][28] ) );
  DFFARX1 \FIFO_reg[42][27]  ( .D(n3214), .CLK(clk_in), .RSTB(n7181), .Q(
        \FIFO[42][27] ) );
  DFFARX1 \FIFO_reg[42][26]  ( .D(n3213), .CLK(clk_in), .RSTB(n7181), .Q(
        \FIFO[42][26] ) );
  DFFARX1 \FIFO_reg[42][25]  ( .D(n3212), .CLK(clk_in), .RSTB(n7181), .Q(
        \FIFO[42][25] ) );
  DFFARX1 \FIFO_reg[42][24]  ( .D(n3211), .CLK(clk_in), .RSTB(n7181), .Q(
        \FIFO[42][24] ) );
  DFFARX1 \FIFO_reg[42][23]  ( .D(n3210), .CLK(clk_in), .RSTB(n7181), .Q(
        \FIFO[42][23] ) );
  DFFARX1 \FIFO_reg[42][22]  ( .D(n3209), .CLK(clk_in), .RSTB(n7181), .Q(
        \FIFO[42][22] ) );
  DFFARX1 \FIFO_reg[42][21]  ( .D(n3208), .CLK(clk_in), .RSTB(n7181), .Q(
        \FIFO[42][21] ) );
  DFFARX1 \FIFO_reg[42][20]  ( .D(n3207), .CLK(clk_in), .RSTB(n7181), .Q(
        \FIFO[42][20] ) );
  DFFARX1 \FIFO_reg[42][19]  ( .D(n3206), .CLK(clk_in), .RSTB(n7182), .Q(
        \FIFO[42][19] ) );
  DFFARX1 \FIFO_reg[42][18]  ( .D(n3205), .CLK(clk_in), .RSTB(n7182), .Q(
        \FIFO[42][18] ) );
  DFFARX1 \FIFO_reg[42][17]  ( .D(n3204), .CLK(clk_in), .RSTB(n7182), .Q(
        \FIFO[42][17] ) );
  DFFARX1 \FIFO_reg[42][16]  ( .D(n3203), .CLK(clk_in), .RSTB(n7182), .Q(
        \FIFO[42][16] ) );
  DFFARX1 \FIFO_reg[42][15]  ( .D(n3202), .CLK(clk_in), .RSTB(n7182), .Q(
        \FIFO[42][15] ) );
  DFFARX1 \FIFO_reg[42][14]  ( .D(n3201), .CLK(clk_in), .RSTB(n7182), .Q(
        \FIFO[42][14] ) );
  DFFARX1 \FIFO_reg[42][13]  ( .D(n3200), .CLK(clk_in), .RSTB(n7182), .Q(
        \FIFO[42][13] ) );
  DFFARX1 \FIFO_reg[42][12]  ( .D(n3199), .CLK(clk_in), .RSTB(n7182), .Q(
        \FIFO[42][12] ) );
  DFFARX1 \FIFO_reg[42][11]  ( .D(n3198), .CLK(clk_in), .RSTB(n7182), .Q(
        \FIFO[42][11] ) );
  DFFARX1 \FIFO_reg[42][10]  ( .D(n3197), .CLK(clk_in), .RSTB(n7182), .Q(
        \FIFO[42][10] ) );
  DFFARX1 \FIFO_reg[42][9]  ( .D(n3196), .CLK(clk_in), .RSTB(n7182), .Q(
        \FIFO[42][9] ) );
  DFFARX1 \FIFO_reg[42][8]  ( .D(n3195), .CLK(clk_in), .RSTB(n7182), .Q(
        \FIFO[42][8] ) );
  DFFARX1 \FIFO_reg[42][7]  ( .D(n3194), .CLK(clk_in), .RSTB(n7182), .Q(
        \FIFO[42][7] ) );
  DFFARX1 \FIFO_reg[42][6]  ( .D(n3193), .CLK(clk_in), .RSTB(n7182), .Q(
        \FIFO[42][6] ) );
  DFFARX1 \FIFO_reg[42][5]  ( .D(n3192), .CLK(clk_in), .RSTB(n7182), .Q(
        \FIFO[42][5] ) );
  DFFARX1 \FIFO_reg[42][4]  ( .D(n3191), .CLK(clk_in), .RSTB(n7182), .Q(
        \FIFO[42][4] ) );
  DFFARX1 \FIFO_reg[42][3]  ( .D(n3190), .CLK(clk_in), .RSTB(n7182), .Q(
        \FIFO[42][3] ) );
  DFFARX1 \FIFO_reg[42][2]  ( .D(n3189), .CLK(clk_in), .RSTB(n7182), .Q(
        \FIFO[42][2] ) );
  DFFARX1 \FIFO_reg[42][1]  ( .D(n3188), .CLK(clk_in), .RSTB(n7183), .Q(
        \FIFO[42][1] ) );
  DFFARX1 \FIFO_reg[42][0]  ( .D(n3187), .CLK(clk_in), .RSTB(n7183), .Q(
        \FIFO[42][0] ) );
  DFFARX1 \FIFO_reg[43][31]  ( .D(n3186), .CLK(clk_in), .RSTB(n7183), .Q(
        \FIFO[43][31] ) );
  DFFARX1 \FIFO_reg[43][30]  ( .D(n3185), .CLK(clk_in), .RSTB(n7183), .Q(
        \FIFO[43][30] ) );
  DFFARX1 \FIFO_reg[43][29]  ( .D(n3184), .CLK(clk_in), .RSTB(n7183), .Q(
        \FIFO[43][29] ) );
  DFFARX1 \FIFO_reg[43][28]  ( .D(n3183), .CLK(clk_in), .RSTB(n7183), .Q(
        \FIFO[43][28] ) );
  DFFARX1 \FIFO_reg[43][27]  ( .D(n3182), .CLK(clk_in), .RSTB(n7183), .Q(
        \FIFO[43][27] ) );
  DFFARX1 \FIFO_reg[43][26]  ( .D(n3181), .CLK(clk_in), .RSTB(n7183), .Q(
        \FIFO[43][26] ) );
  DFFARX1 \FIFO_reg[43][25]  ( .D(n3180), .CLK(clk_in), .RSTB(n7183), .Q(
        \FIFO[43][25] ) );
  DFFARX1 \FIFO_reg[43][24]  ( .D(n3179), .CLK(clk_in), .RSTB(n7183), .Q(
        \FIFO[43][24] ) );
  DFFARX1 \FIFO_reg[43][23]  ( .D(n3178), .CLK(clk_in), .RSTB(n7183), .Q(
        \FIFO[43][23] ) );
  DFFARX1 \FIFO_reg[43][22]  ( .D(n3177), .CLK(clk_in), .RSTB(n7183), .Q(
        \FIFO[43][22] ) );
  DFFARX1 \FIFO_reg[43][21]  ( .D(n3176), .CLK(clk_in), .RSTB(n7183), .Q(
        \FIFO[43][21] ) );
  DFFARX1 \FIFO_reg[43][20]  ( .D(n3175), .CLK(clk_in), .RSTB(n7183), .Q(
        \FIFO[43][20] ) );
  DFFARX1 \FIFO_reg[43][19]  ( .D(n3174), .CLK(clk_in), .RSTB(n7183), .Q(
        \FIFO[43][19] ) );
  DFFARX1 \FIFO_reg[43][18]  ( .D(n3173), .CLK(clk_in), .RSTB(n7183), .Q(
        \FIFO[43][18] ) );
  DFFARX1 \FIFO_reg[43][17]  ( .D(n3172), .CLK(clk_in), .RSTB(n7183), .Q(
        \FIFO[43][17] ) );
  DFFARX1 \FIFO_reg[43][16]  ( .D(n3171), .CLK(clk_in), .RSTB(n7183), .Q(
        \FIFO[43][16] ) );
  DFFARX1 \FIFO_reg[43][15]  ( .D(n3170), .CLK(clk_in), .RSTB(n7184), .Q(
        \FIFO[43][15] ) );
  DFFARX1 \FIFO_reg[43][14]  ( .D(n3169), .CLK(clk_in), .RSTB(n7184), .Q(
        \FIFO[43][14] ) );
  DFFARX1 \FIFO_reg[43][13]  ( .D(n3168), .CLK(clk_in), .RSTB(n7184), .Q(
        \FIFO[43][13] ) );
  DFFARX1 \FIFO_reg[43][12]  ( .D(n3167), .CLK(clk_in), .RSTB(n7184), .Q(
        \FIFO[43][12] ) );
  DFFARX1 \FIFO_reg[43][11]  ( .D(n3166), .CLK(clk_in), .RSTB(n7184), .Q(
        \FIFO[43][11] ) );
  DFFARX1 \FIFO_reg[43][10]  ( .D(n3165), .CLK(clk_in), .RSTB(n7184), .Q(
        \FIFO[43][10] ) );
  DFFARX1 \FIFO_reg[43][9]  ( .D(n3164), .CLK(clk_in), .RSTB(n7184), .Q(
        \FIFO[43][9] ) );
  DFFARX1 \FIFO_reg[43][8]  ( .D(n3163), .CLK(clk_in), .RSTB(n7184), .Q(
        \FIFO[43][8] ) );
  DFFARX1 \FIFO_reg[43][7]  ( .D(n3162), .CLK(clk_in), .RSTB(n7184), .Q(
        \FIFO[43][7] ) );
  DFFARX1 \FIFO_reg[43][6]  ( .D(n3161), .CLK(clk_in), .RSTB(n7184), .Q(
        \FIFO[43][6] ) );
  DFFARX1 \FIFO_reg[43][5]  ( .D(n3160), .CLK(clk_in), .RSTB(n7184), .Q(
        \FIFO[43][5] ) );
  DFFARX1 \FIFO_reg[43][4]  ( .D(n3159), .CLK(clk_in), .RSTB(n7184), .Q(
        \FIFO[43][4] ) );
  DFFARX1 \FIFO_reg[43][3]  ( .D(n3158), .CLK(clk_in), .RSTB(n7184), .Q(
        \FIFO[43][3] ) );
  DFFARX1 \FIFO_reg[43][2]  ( .D(n3157), .CLK(clk_in), .RSTB(n7184), .Q(
        \FIFO[43][2] ) );
  DFFARX1 \FIFO_reg[43][1]  ( .D(n3156), .CLK(clk_in), .RSTB(n7184), .Q(
        \FIFO[43][1] ) );
  DFFARX1 \FIFO_reg[43][0]  ( .D(n3155), .CLK(clk_in), .RSTB(n7184), .Q(
        \FIFO[43][0] ) );
  DFFARX1 \FIFO_reg[44][31]  ( .D(n3154), .CLK(clk_in), .RSTB(n7184), .Q(
        \FIFO[44][31] ) );
  DFFARX1 \FIFO_reg[44][30]  ( .D(n3153), .CLK(clk_in), .RSTB(n7184), .Q(
        \FIFO[44][30] ) );
  DFFARX1 \FIFO_reg[44][29]  ( .D(n3152), .CLK(clk_in), .RSTB(n7185), .Q(
        \FIFO[44][29] ) );
  DFFARX1 \FIFO_reg[44][28]  ( .D(n3151), .CLK(clk_in), .RSTB(n7185), .Q(
        \FIFO[44][28] ) );
  DFFARX1 \FIFO_reg[44][27]  ( .D(n3150), .CLK(clk_in), .RSTB(n7185), .Q(
        \FIFO[44][27] ) );
  DFFARX1 \FIFO_reg[44][26]  ( .D(n3149), .CLK(clk_in), .RSTB(n7185), .Q(
        \FIFO[44][26] ) );
  DFFARX1 \FIFO_reg[44][25]  ( .D(n3148), .CLK(clk_in), .RSTB(n7185), .Q(
        \FIFO[44][25] ) );
  DFFARX1 \FIFO_reg[44][24]  ( .D(n3147), .CLK(clk_in), .RSTB(n7185), .Q(
        \FIFO[44][24] ) );
  DFFARX1 \FIFO_reg[44][23]  ( .D(n3146), .CLK(clk_in), .RSTB(n7185), .Q(
        \FIFO[44][23] ) );
  DFFARX1 \FIFO_reg[44][22]  ( .D(n3145), .CLK(clk_in), .RSTB(n7185), .Q(
        \FIFO[44][22] ) );
  DFFARX1 \FIFO_reg[44][21]  ( .D(n3144), .CLK(clk_in), .RSTB(n7185), .Q(
        \FIFO[44][21] ) );
  DFFARX1 \FIFO_reg[44][20]  ( .D(n3143), .CLK(clk_in), .RSTB(n7185), .Q(
        \FIFO[44][20] ) );
  DFFARX1 \FIFO_reg[44][19]  ( .D(n3142), .CLK(clk_in), .RSTB(n7185), .Q(
        \FIFO[44][19] ) );
  DFFARX1 \FIFO_reg[44][18]  ( .D(n3141), .CLK(clk_in), .RSTB(n7185), .Q(
        \FIFO[44][18] ) );
  DFFARX1 \FIFO_reg[44][17]  ( .D(n3140), .CLK(clk_in), .RSTB(n7185), .Q(
        \FIFO[44][17] ) );
  DFFARX1 \FIFO_reg[44][16]  ( .D(n3139), .CLK(clk_in), .RSTB(n7185), .Q(
        \FIFO[44][16] ) );
  DFFARX1 \FIFO_reg[44][15]  ( .D(n3138), .CLK(clk_in), .RSTB(n7185), .Q(
        \FIFO[44][15] ) );
  DFFARX1 \FIFO_reg[44][14]  ( .D(n3137), .CLK(clk_in), .RSTB(n7185), .Q(
        \FIFO[44][14] ) );
  DFFARX1 \FIFO_reg[44][13]  ( .D(n3136), .CLK(clk_in), .RSTB(n7185), .Q(
        \FIFO[44][13] ) );
  DFFARX1 \FIFO_reg[44][12]  ( .D(n3135), .CLK(clk_in), .RSTB(n7185), .Q(
        \FIFO[44][12] ) );
  DFFARX1 \FIFO_reg[44][11]  ( .D(n3134), .CLK(clk_in), .RSTB(n7186), .Q(
        \FIFO[44][11] ) );
  DFFARX1 \FIFO_reg[44][10]  ( .D(n3133), .CLK(clk_in), .RSTB(n7186), .Q(
        \FIFO[44][10] ) );
  DFFARX1 \FIFO_reg[44][9]  ( .D(n3132), .CLK(clk_in), .RSTB(n7186), .Q(
        \FIFO[44][9] ) );
  DFFARX1 \FIFO_reg[44][8]  ( .D(n3131), .CLK(clk_in), .RSTB(n7186), .Q(
        \FIFO[44][8] ) );
  DFFARX1 \FIFO_reg[44][7]  ( .D(n3130), .CLK(clk_in), .RSTB(n7186), .Q(
        \FIFO[44][7] ) );
  DFFARX1 \FIFO_reg[44][6]  ( .D(n3129), .CLK(clk_in), .RSTB(n7186), .Q(
        \FIFO[44][6] ) );
  DFFARX1 \FIFO_reg[44][5]  ( .D(n3128), .CLK(clk_in), .RSTB(n7186), .Q(
        \FIFO[44][5] ) );
  DFFARX1 \FIFO_reg[44][4]  ( .D(n3127), .CLK(clk_in), .RSTB(n7186), .Q(
        \FIFO[44][4] ) );
  DFFARX1 \FIFO_reg[44][3]  ( .D(n3126), .CLK(clk_in), .RSTB(n7186), .Q(
        \FIFO[44][3] ) );
  DFFARX1 \FIFO_reg[44][2]  ( .D(n3125), .CLK(clk_in), .RSTB(n7186), .Q(
        \FIFO[44][2] ) );
  DFFARX1 \FIFO_reg[44][1]  ( .D(n3124), .CLK(clk_in), .RSTB(n7186), .Q(
        \FIFO[44][1] ) );
  DFFARX1 \FIFO_reg[44][0]  ( .D(n3123), .CLK(clk_in), .RSTB(n7186), .Q(
        \FIFO[44][0] ) );
  DFFARX1 \FIFO_reg[45][31]  ( .D(n3122), .CLK(clk_in), .RSTB(n7186), .Q(
        \FIFO[45][31] ) );
  DFFARX1 \FIFO_reg[45][30]  ( .D(n3121), .CLK(clk_in), .RSTB(n7186), .Q(
        \FIFO[45][30] ) );
  DFFARX1 \FIFO_reg[45][29]  ( .D(n3120), .CLK(clk_in), .RSTB(n7186), .Q(
        \FIFO[45][29] ) );
  DFFARX1 \FIFO_reg[45][28]  ( .D(n3119), .CLK(clk_in), .RSTB(n7186), .Q(
        \FIFO[45][28] ) );
  DFFARX1 \FIFO_reg[45][27]  ( .D(n3118), .CLK(clk_in), .RSTB(n7186), .Q(
        \FIFO[45][27] ) );
  DFFARX1 \FIFO_reg[45][26]  ( .D(n3117), .CLK(clk_in), .RSTB(n7186), .Q(
        \FIFO[45][26] ) );
  DFFARX1 \FIFO_reg[45][25]  ( .D(n3116), .CLK(clk_in), .RSTB(n7187), .Q(
        \FIFO[45][25] ) );
  DFFARX1 \FIFO_reg[45][24]  ( .D(n3115), .CLK(clk_in), .RSTB(n7187), .Q(
        \FIFO[45][24] ) );
  DFFARX1 \FIFO_reg[45][23]  ( .D(n3114), .CLK(clk_in), .RSTB(n7187), .Q(
        \FIFO[45][23] ) );
  DFFARX1 \FIFO_reg[45][22]  ( .D(n3113), .CLK(clk_in), .RSTB(n7187), .Q(
        \FIFO[45][22] ) );
  DFFARX1 \FIFO_reg[45][21]  ( .D(n3112), .CLK(clk_in), .RSTB(n7187), .Q(
        \FIFO[45][21] ) );
  DFFARX1 \FIFO_reg[45][20]  ( .D(n3111), .CLK(clk_in), .RSTB(n7187), .Q(
        \FIFO[45][20] ) );
  DFFARX1 \FIFO_reg[45][19]  ( .D(n3110), .CLK(clk_in), .RSTB(n7187), .Q(
        \FIFO[45][19] ) );
  DFFARX1 \FIFO_reg[45][18]  ( .D(n3109), .CLK(clk_in), .RSTB(n7187), .Q(
        \FIFO[45][18] ) );
  DFFARX1 \FIFO_reg[45][17]  ( .D(n3108), .CLK(clk_in), .RSTB(n7187), .Q(
        \FIFO[45][17] ) );
  DFFARX1 \FIFO_reg[45][16]  ( .D(n3107), .CLK(clk_in), .RSTB(n7187), .Q(
        \FIFO[45][16] ) );
  DFFARX1 \FIFO_reg[45][15]  ( .D(n3106), .CLK(clk_in), .RSTB(n7187), .Q(
        \FIFO[45][15] ) );
  DFFARX1 \FIFO_reg[45][14]  ( .D(n3105), .CLK(clk_in), .RSTB(n7187), .Q(
        \FIFO[45][14] ) );
  DFFARX1 \FIFO_reg[45][13]  ( .D(n3104), .CLK(clk_in), .RSTB(n7187), .Q(
        \FIFO[45][13] ) );
  DFFARX1 \FIFO_reg[45][12]  ( .D(n3103), .CLK(clk_in), .RSTB(n7187), .Q(
        \FIFO[45][12] ) );
  DFFARX1 \FIFO_reg[45][11]  ( .D(n3102), .CLK(clk_in), .RSTB(n7187), .Q(
        \FIFO[45][11] ) );
  DFFARX1 \FIFO_reg[45][10]  ( .D(n3101), .CLK(clk_in), .RSTB(n7187), .Q(
        \FIFO[45][10] ) );
  DFFARX1 \FIFO_reg[45][9]  ( .D(n3100), .CLK(clk_in), .RSTB(n7187), .Q(
        \FIFO[45][9] ) );
  DFFARX1 \FIFO_reg[45][8]  ( .D(n3099), .CLK(clk_in), .RSTB(n7187), .Q(
        \FIFO[45][8] ) );
  DFFARX1 \FIFO_reg[45][7]  ( .D(n3098), .CLK(clk_in), .RSTB(n7188), .Q(
        \FIFO[45][7] ) );
  DFFARX1 \FIFO_reg[45][6]  ( .D(n3097), .CLK(clk_in), .RSTB(n7188), .Q(
        \FIFO[45][6] ) );
  DFFARX1 \FIFO_reg[45][5]  ( .D(n3096), .CLK(clk_in), .RSTB(n7188), .Q(
        \FIFO[45][5] ) );
  DFFARX1 \FIFO_reg[45][4]  ( .D(n3095), .CLK(clk_in), .RSTB(n7188), .Q(
        \FIFO[45][4] ) );
  DFFARX1 \FIFO_reg[45][3]  ( .D(n3094), .CLK(clk_in), .RSTB(n7188), .Q(
        \FIFO[45][3] ) );
  DFFARX1 \FIFO_reg[45][2]  ( .D(n3093), .CLK(clk_in), .RSTB(n7188), .Q(
        \FIFO[45][2] ) );
  DFFARX1 \FIFO_reg[45][1]  ( .D(n3092), .CLK(clk_in), .RSTB(n7188), .Q(
        \FIFO[45][1] ) );
  DFFARX1 \FIFO_reg[45][0]  ( .D(n3091), .CLK(clk_in), .RSTB(n7188), .Q(
        \FIFO[45][0] ) );
  DFFARX1 \FIFO_reg[46][31]  ( .D(n3090), .CLK(clk_in), .RSTB(n7188), .Q(
        \FIFO[46][31] ) );
  DFFARX1 \FIFO_reg[46][30]  ( .D(n3089), .CLK(clk_in), .RSTB(n7188), .Q(
        \FIFO[46][30] ) );
  DFFARX1 \FIFO_reg[46][29]  ( .D(n3088), .CLK(clk_in), .RSTB(n7188), .Q(
        \FIFO[46][29] ) );
  DFFARX1 \FIFO_reg[46][28]  ( .D(n3087), .CLK(clk_in), .RSTB(n7188), .Q(
        \FIFO[46][28] ) );
  DFFARX1 \FIFO_reg[46][27]  ( .D(n3086), .CLK(clk_in), .RSTB(n7188), .Q(
        \FIFO[46][27] ) );
  DFFARX1 \FIFO_reg[46][26]  ( .D(n3085), .CLK(clk_in), .RSTB(n7188), .Q(
        \FIFO[46][26] ) );
  DFFARX1 \FIFO_reg[46][25]  ( .D(n3084), .CLK(clk_in), .RSTB(n7188), .Q(
        \FIFO[46][25] ) );
  DFFARX1 \FIFO_reg[46][24]  ( .D(n3083), .CLK(clk_in), .RSTB(n7188), .Q(
        \FIFO[46][24] ) );
  DFFARX1 \FIFO_reg[46][23]  ( .D(n3082), .CLK(clk_in), .RSTB(n7188), .Q(
        \FIFO[46][23] ) );
  DFFARX1 \FIFO_reg[46][22]  ( .D(n3081), .CLK(clk_in), .RSTB(n7188), .Q(
        \FIFO[46][22] ) );
  DFFARX1 \FIFO_reg[46][21]  ( .D(n3080), .CLK(clk_in), .RSTB(n7189), .Q(
        \FIFO[46][21] ) );
  DFFARX1 \FIFO_reg[46][20]  ( .D(n3079), .CLK(clk_in), .RSTB(n7189), .Q(
        \FIFO[46][20] ) );
  DFFARX1 \FIFO_reg[46][19]  ( .D(n3078), .CLK(clk_in), .RSTB(n7189), .Q(
        \FIFO[46][19] ) );
  DFFARX1 \FIFO_reg[46][18]  ( .D(n3077), .CLK(clk_in), .RSTB(n7189), .Q(
        \FIFO[46][18] ) );
  DFFARX1 \FIFO_reg[46][17]  ( .D(n3076), .CLK(clk_in), .RSTB(n7189), .Q(
        \FIFO[46][17] ) );
  DFFARX1 \FIFO_reg[46][16]  ( .D(n3075), .CLK(clk_in), .RSTB(n7189), .Q(
        \FIFO[46][16] ) );
  DFFARX1 \FIFO_reg[46][15]  ( .D(n3074), .CLK(clk_in), .RSTB(n7189), .Q(
        \FIFO[46][15] ) );
  DFFARX1 \FIFO_reg[46][14]  ( .D(n3073), .CLK(clk_in), .RSTB(n7189), .Q(
        \FIFO[46][14] ) );
  DFFARX1 \FIFO_reg[46][13]  ( .D(n3072), .CLK(clk_in), .RSTB(n7189), .Q(
        \FIFO[46][13] ) );
  DFFARX1 \FIFO_reg[46][12]  ( .D(n3071), .CLK(clk_in), .RSTB(n7189), .Q(
        \FIFO[46][12] ) );
  DFFARX1 \FIFO_reg[46][11]  ( .D(n3070), .CLK(clk_in), .RSTB(n7189), .Q(
        \FIFO[46][11] ) );
  DFFARX1 \FIFO_reg[46][10]  ( .D(n3069), .CLK(clk_in), .RSTB(n7189), .Q(
        \FIFO[46][10] ) );
  DFFARX1 \FIFO_reg[46][9]  ( .D(n3068), .CLK(clk_in), .RSTB(n7189), .Q(
        \FIFO[46][9] ) );
  DFFARX1 \FIFO_reg[46][8]  ( .D(n3067), .CLK(clk_in), .RSTB(n7189), .Q(
        \FIFO[46][8] ) );
  DFFARX1 \FIFO_reg[46][7]  ( .D(n3066), .CLK(clk_in), .RSTB(n7189), .Q(
        \FIFO[46][7] ) );
  DFFARX1 \FIFO_reg[46][6]  ( .D(n3065), .CLK(clk_in), .RSTB(n7189), .Q(
        \FIFO[46][6] ) );
  DFFARX1 \FIFO_reg[46][5]  ( .D(n3064), .CLK(clk_in), .RSTB(n7189), .Q(
        \FIFO[46][5] ) );
  DFFARX1 \FIFO_reg[46][4]  ( .D(n3063), .CLK(clk_in), .RSTB(n7189), .Q(
        \FIFO[46][4] ) );
  DFFARX1 \FIFO_reg[46][3]  ( .D(n3062), .CLK(clk_in), .RSTB(n7190), .Q(
        \FIFO[46][3] ) );
  DFFARX1 \FIFO_reg[46][2]  ( .D(n3061), .CLK(clk_in), .RSTB(n7190), .Q(
        \FIFO[46][2] ) );
  DFFARX1 \FIFO_reg[46][1]  ( .D(n3060), .CLK(clk_in), .RSTB(n7190), .Q(
        \FIFO[46][1] ) );
  DFFARX1 \FIFO_reg[46][0]  ( .D(n3059), .CLK(clk_in), .RSTB(n7190), .Q(
        \FIFO[46][0] ) );
  DFFARX1 \FIFO_reg[47][31]  ( .D(n3058), .CLK(clk_in), .RSTB(n7190), .Q(
        \FIFO[47][31] ) );
  DFFARX1 \FIFO_reg[47][30]  ( .D(n3057), .CLK(clk_in), .RSTB(n7190), .Q(
        \FIFO[47][30] ) );
  DFFARX1 \FIFO_reg[47][29]  ( .D(n3056), .CLK(clk_in), .RSTB(n7190), .Q(
        \FIFO[47][29] ) );
  DFFARX1 \FIFO_reg[47][28]  ( .D(n3055), .CLK(clk_in), .RSTB(n7190), .Q(
        \FIFO[47][28] ) );
  DFFARX1 \FIFO_reg[47][27]  ( .D(n3054), .CLK(clk_in), .RSTB(n7190), .Q(
        \FIFO[47][27] ) );
  DFFARX1 \FIFO_reg[47][26]  ( .D(n3053), .CLK(clk_in), .RSTB(n7190), .Q(
        \FIFO[47][26] ) );
  DFFARX1 \FIFO_reg[47][25]  ( .D(n3052), .CLK(clk_in), .RSTB(n7190), .Q(
        \FIFO[47][25] ) );
  DFFARX1 \FIFO_reg[47][24]  ( .D(n3051), .CLK(clk_in), .RSTB(n7190), .Q(
        \FIFO[47][24] ) );
  DFFARX1 \FIFO_reg[47][23]  ( .D(n3050), .CLK(clk_in), .RSTB(n7190), .Q(
        \FIFO[47][23] ) );
  DFFARX1 \FIFO_reg[47][22]  ( .D(n3049), .CLK(clk_in), .RSTB(n7190), .Q(
        \FIFO[47][22] ) );
  DFFARX1 \FIFO_reg[47][21]  ( .D(n3048), .CLK(clk_in), .RSTB(n7190), .Q(
        \FIFO[47][21] ) );
  DFFARX1 \FIFO_reg[47][20]  ( .D(n3047), .CLK(clk_in), .RSTB(n7190), .Q(
        \FIFO[47][20] ) );
  DFFARX1 \FIFO_reg[47][19]  ( .D(n3046), .CLK(clk_in), .RSTB(n7190), .Q(
        \FIFO[47][19] ) );
  DFFARX1 \FIFO_reg[47][18]  ( .D(n3045), .CLK(clk_in), .RSTB(n7190), .Q(
        \FIFO[47][18] ) );
  DFFARX1 \FIFO_reg[47][17]  ( .D(n3044), .CLK(clk_in), .RSTB(n7191), .Q(
        \FIFO[47][17] ) );
  DFFARX1 \FIFO_reg[47][16]  ( .D(n3043), .CLK(clk_in), .RSTB(n7191), .Q(
        \FIFO[47][16] ) );
  DFFARX1 \FIFO_reg[47][15]  ( .D(n3042), .CLK(clk_in), .RSTB(n7191), .Q(
        \FIFO[47][15] ) );
  DFFARX1 \FIFO_reg[47][14]  ( .D(n3041), .CLK(clk_in), .RSTB(n7191), .Q(
        \FIFO[47][14] ) );
  DFFARX1 \FIFO_reg[47][13]  ( .D(n3040), .CLK(clk_in), .RSTB(n7191), .Q(
        \FIFO[47][13] ) );
  DFFARX1 \FIFO_reg[47][12]  ( .D(n3039), .CLK(clk_in), .RSTB(n7191), .Q(
        \FIFO[47][12] ) );
  DFFARX1 \FIFO_reg[47][11]  ( .D(n3038), .CLK(clk_in), .RSTB(n7191), .Q(
        \FIFO[47][11] ) );
  DFFARX1 \FIFO_reg[47][10]  ( .D(n3037), .CLK(clk_in), .RSTB(n7191), .Q(
        \FIFO[47][10] ) );
  DFFARX1 \FIFO_reg[47][9]  ( .D(n3036), .CLK(clk_in), .RSTB(n7191), .Q(
        \FIFO[47][9] ) );
  DFFARX1 \FIFO_reg[47][8]  ( .D(n3035), .CLK(clk_in), .RSTB(n7191), .Q(
        \FIFO[47][8] ) );
  DFFARX1 \FIFO_reg[47][7]  ( .D(n3034), .CLK(clk_in), .RSTB(n7191), .Q(
        \FIFO[47][7] ) );
  DFFARX1 \FIFO_reg[47][6]  ( .D(n3033), .CLK(clk_in), .RSTB(n7191), .Q(
        \FIFO[47][6] ) );
  DFFARX1 \FIFO_reg[47][5]  ( .D(n3032), .CLK(clk_in), .RSTB(n7191), .Q(
        \FIFO[47][5] ) );
  DFFARX1 \FIFO_reg[47][4]  ( .D(n3031), .CLK(clk_in), .RSTB(n7191), .Q(
        \FIFO[47][4] ) );
  DFFARX1 \FIFO_reg[47][3]  ( .D(n3030), .CLK(clk_in), .RSTB(n7191), .Q(
        \FIFO[47][3] ) );
  DFFARX1 \FIFO_reg[47][2]  ( .D(n3029), .CLK(clk_in), .RSTB(n7191), .Q(
        \FIFO[47][2] ) );
  DFFARX1 \FIFO_reg[47][1]  ( .D(n3028), .CLK(clk_in), .RSTB(n7191), .Q(
        \FIFO[47][1] ) );
  DFFARX1 \FIFO_reg[47][0]  ( .D(n3027), .CLK(clk_in), .RSTB(n7191), .Q(
        \FIFO[47][0] ) );
  DFFARX1 \FIFO_reg[48][31]  ( .D(n3026), .CLK(clk_in), .RSTB(n7192), .Q(
        \FIFO[48][31] ) );
  DFFARX1 \FIFO_reg[48][30]  ( .D(n3025), .CLK(clk_in), .RSTB(n7192), .Q(
        \FIFO[48][30] ) );
  DFFARX1 \FIFO_reg[48][29]  ( .D(n3024), .CLK(clk_in), .RSTB(n7192), .Q(
        \FIFO[48][29] ) );
  DFFARX1 \FIFO_reg[48][28]  ( .D(n3023), .CLK(clk_in), .RSTB(n7192), .Q(
        \FIFO[48][28] ) );
  DFFARX1 \FIFO_reg[48][27]  ( .D(n3022), .CLK(clk_in), .RSTB(n7192), .Q(
        \FIFO[48][27] ) );
  DFFARX1 \FIFO_reg[48][26]  ( .D(n3021), .CLK(clk_in), .RSTB(n7192), .Q(
        \FIFO[48][26] ) );
  DFFARX1 \FIFO_reg[48][25]  ( .D(n3020), .CLK(clk_in), .RSTB(n7192), .Q(
        \FIFO[48][25] ) );
  DFFARX1 \FIFO_reg[48][24]  ( .D(n3019), .CLK(clk_in), .RSTB(n7192), .Q(
        \FIFO[48][24] ) );
  DFFARX1 \FIFO_reg[48][23]  ( .D(n3018), .CLK(clk_in), .RSTB(n7192), .Q(
        \FIFO[48][23] ) );
  DFFARX1 \FIFO_reg[48][22]  ( .D(n3017), .CLK(clk_in), .RSTB(n7192), .Q(
        \FIFO[48][22] ) );
  DFFARX1 \FIFO_reg[48][21]  ( .D(n3016), .CLK(clk_in), .RSTB(n7192), .Q(
        \FIFO[48][21] ) );
  DFFARX1 \FIFO_reg[48][20]  ( .D(n3015), .CLK(clk_in), .RSTB(n7192), .Q(
        \FIFO[48][20] ) );
  DFFARX1 \FIFO_reg[48][19]  ( .D(n3014), .CLK(clk_in), .RSTB(n7192), .Q(
        \FIFO[48][19] ) );
  DFFARX1 \FIFO_reg[48][18]  ( .D(n3013), .CLK(clk_in), .RSTB(n7192), .Q(
        \FIFO[48][18] ) );
  DFFARX1 \FIFO_reg[48][17]  ( .D(n3012), .CLK(clk_in), .RSTB(n7192), .Q(
        \FIFO[48][17] ) );
  DFFARX1 \FIFO_reg[48][16]  ( .D(n3011), .CLK(clk_in), .RSTB(n7192), .Q(
        \FIFO[48][16] ) );
  DFFARX1 \FIFO_reg[48][15]  ( .D(n3010), .CLK(clk_in), .RSTB(n7192), .Q(
        \FIFO[48][15] ) );
  DFFARX1 \FIFO_reg[48][14]  ( .D(n3009), .CLK(clk_in), .RSTB(n7192), .Q(
        \FIFO[48][14] ) );
  DFFARX1 \FIFO_reg[48][13]  ( .D(n3008), .CLK(clk_in), .RSTB(n7193), .Q(
        \FIFO[48][13] ) );
  DFFARX1 \FIFO_reg[48][12]  ( .D(n3007), .CLK(clk_in), .RSTB(n7193), .Q(
        \FIFO[48][12] ) );
  DFFARX1 \FIFO_reg[48][11]  ( .D(n3006), .CLK(clk_in), .RSTB(n7193), .Q(
        \FIFO[48][11] ) );
  DFFARX1 \FIFO_reg[48][10]  ( .D(n3005), .CLK(clk_in), .RSTB(n7193), .Q(
        \FIFO[48][10] ) );
  DFFARX1 \FIFO_reg[48][9]  ( .D(n3004), .CLK(clk_in), .RSTB(n7193), .Q(
        \FIFO[48][9] ) );
  DFFARX1 \FIFO_reg[48][8]  ( .D(n3003), .CLK(clk_in), .RSTB(n7193), .Q(
        \FIFO[48][8] ) );
  DFFARX1 \FIFO_reg[48][7]  ( .D(n3002), .CLK(clk_in), .RSTB(n7193), .Q(
        \FIFO[48][7] ) );
  DFFARX1 \FIFO_reg[48][6]  ( .D(n3001), .CLK(clk_in), .RSTB(n7193), .Q(
        \FIFO[48][6] ) );
  DFFARX1 \FIFO_reg[48][5]  ( .D(n3000), .CLK(clk_in), .RSTB(n7193), .Q(
        \FIFO[48][5] ) );
  DFFARX1 \FIFO_reg[48][4]  ( .D(n2999), .CLK(clk_in), .RSTB(n7193), .Q(
        \FIFO[48][4] ) );
  DFFARX1 \FIFO_reg[48][3]  ( .D(n2998), .CLK(clk_in), .RSTB(n7193), .Q(
        \FIFO[48][3] ) );
  DFFARX1 \FIFO_reg[48][2]  ( .D(n2997), .CLK(clk_in), .RSTB(n7193), .Q(
        \FIFO[48][2] ) );
  DFFARX1 \FIFO_reg[48][1]  ( .D(n2996), .CLK(clk_in), .RSTB(n7193), .Q(
        \FIFO[48][1] ) );
  DFFARX1 \FIFO_reg[48][0]  ( .D(n2995), .CLK(clk_in), .RSTB(n7193), .Q(
        \FIFO[48][0] ) );
  DFFARX1 \FIFO_reg[49][31]  ( .D(n2994), .CLK(clk_in), .RSTB(n7193), .Q(
        \FIFO[49][31] ) );
  DFFARX1 \FIFO_reg[49][30]  ( .D(n2993), .CLK(clk_in), .RSTB(n7193), .Q(
        \FIFO[49][30] ) );
  DFFARX1 \FIFO_reg[49][29]  ( .D(n2992), .CLK(clk_in), .RSTB(n7193), .Q(
        \FIFO[49][29] ) );
  DFFARX1 \FIFO_reg[49][28]  ( .D(n2991), .CLK(clk_in), .RSTB(n7193), .Q(
        \FIFO[49][28] ) );
  DFFARX1 \FIFO_reg[49][27]  ( .D(n2990), .CLK(clk_in), .RSTB(n7194), .Q(
        \FIFO[49][27] ) );
  DFFARX1 \FIFO_reg[49][26]  ( .D(n2989), .CLK(clk_in), .RSTB(n7194), .Q(
        \FIFO[49][26] ) );
  DFFARX1 \FIFO_reg[49][25]  ( .D(n2988), .CLK(clk_in), .RSTB(n7194), .Q(
        \FIFO[49][25] ) );
  DFFARX1 \FIFO_reg[49][24]  ( .D(n2987), .CLK(clk_in), .RSTB(n7194), .Q(
        \FIFO[49][24] ) );
  DFFARX1 \FIFO_reg[49][23]  ( .D(n2986), .CLK(clk_in), .RSTB(n7194), .Q(
        \FIFO[49][23] ) );
  DFFARX1 \FIFO_reg[49][22]  ( .D(n2985), .CLK(clk_in), .RSTB(n7194), .Q(
        \FIFO[49][22] ) );
  DFFARX1 \FIFO_reg[49][21]  ( .D(n2984), .CLK(clk_in), .RSTB(n7194), .Q(
        \FIFO[49][21] ) );
  DFFARX1 \FIFO_reg[49][20]  ( .D(n2983), .CLK(clk_in), .RSTB(n7194), .Q(
        \FIFO[49][20] ) );
  DFFARX1 \FIFO_reg[49][19]  ( .D(n2982), .CLK(clk_in), .RSTB(n7194), .Q(
        \FIFO[49][19] ) );
  DFFARX1 \FIFO_reg[49][18]  ( .D(n2981), .CLK(clk_in), .RSTB(n7194), .Q(
        \FIFO[49][18] ) );
  DFFARX1 \FIFO_reg[49][17]  ( .D(n2980), .CLK(clk_in), .RSTB(n7194), .Q(
        \FIFO[49][17] ) );
  DFFARX1 \FIFO_reg[49][16]  ( .D(n2979), .CLK(clk_in), .RSTB(n7194), .Q(
        \FIFO[49][16] ) );
  DFFARX1 \FIFO_reg[49][15]  ( .D(n2978), .CLK(clk_in), .RSTB(n7194), .Q(
        \FIFO[49][15] ) );
  DFFARX1 \FIFO_reg[49][14]  ( .D(n2977), .CLK(clk_in), .RSTB(n7194), .Q(
        \FIFO[49][14] ) );
  DFFARX1 \FIFO_reg[49][13]  ( .D(n2976), .CLK(clk_in), .RSTB(n7194), .Q(
        \FIFO[49][13] ) );
  DFFARX1 \FIFO_reg[49][12]  ( .D(n2975), .CLK(clk_in), .RSTB(n7194), .Q(
        \FIFO[49][12] ) );
  DFFARX1 \FIFO_reg[49][11]  ( .D(n2974), .CLK(clk_in), .RSTB(n7194), .Q(
        \FIFO[49][11] ) );
  DFFARX1 \FIFO_reg[49][10]  ( .D(n2973), .CLK(clk_in), .RSTB(n7194), .Q(
        \FIFO[49][10] ) );
  DFFARX1 \FIFO_reg[49][9]  ( .D(n2972), .CLK(clk_in), .RSTB(n7195), .Q(
        \FIFO[49][9] ) );
  DFFARX1 \FIFO_reg[49][8]  ( .D(n2971), .CLK(clk_in), .RSTB(n7195), .Q(
        \FIFO[49][8] ) );
  DFFARX1 \FIFO_reg[49][7]  ( .D(n2970), .CLK(clk_in), .RSTB(n7195), .Q(
        \FIFO[49][7] ) );
  DFFARX1 \FIFO_reg[49][6]  ( .D(n2969), .CLK(clk_in), .RSTB(n7195), .Q(
        \FIFO[49][6] ) );
  DFFARX1 \FIFO_reg[49][5]  ( .D(n2968), .CLK(clk_in), .RSTB(n7195), .Q(
        \FIFO[49][5] ) );
  DFFARX1 \FIFO_reg[49][4]  ( .D(n2967), .CLK(clk_in), .RSTB(n7195), .Q(
        \FIFO[49][4] ) );
  DFFARX1 \FIFO_reg[49][3]  ( .D(n2966), .CLK(clk_in), .RSTB(n7195), .Q(
        \FIFO[49][3] ) );
  DFFARX1 \FIFO_reg[49][2]  ( .D(n2965), .CLK(clk_in), .RSTB(n7195), .Q(
        \FIFO[49][2] ) );
  DFFARX1 \FIFO_reg[49][1]  ( .D(n2964), .CLK(clk_in), .RSTB(n7195), .Q(
        \FIFO[49][1] ) );
  DFFARX1 \FIFO_reg[49][0]  ( .D(n2963), .CLK(clk_in), .RSTB(n7195), .Q(
        \FIFO[49][0] ) );
  DFFARX1 \FIFO_reg[50][31]  ( .D(n2962), .CLK(clk_in), .RSTB(n7195), .Q(
        \FIFO[50][31] ) );
  DFFARX1 \FIFO_reg[50][30]  ( .D(n2961), .CLK(clk_in), .RSTB(n7195), .Q(
        \FIFO[50][30] ) );
  DFFARX1 \FIFO_reg[50][29]  ( .D(n2960), .CLK(clk_in), .RSTB(n7195), .Q(
        \FIFO[50][29] ) );
  DFFARX1 \FIFO_reg[50][28]  ( .D(n2959), .CLK(clk_in), .RSTB(n7195), .Q(
        \FIFO[50][28] ) );
  DFFARX1 \FIFO_reg[50][27]  ( .D(n2958), .CLK(clk_in), .RSTB(n7195), .Q(
        \FIFO[50][27] ) );
  DFFARX1 \FIFO_reg[50][26]  ( .D(n2957), .CLK(clk_in), .RSTB(n7195), .Q(
        \FIFO[50][26] ) );
  DFFARX1 \FIFO_reg[50][25]  ( .D(n2956), .CLK(clk_in), .RSTB(n7195), .Q(
        \FIFO[50][25] ) );
  DFFARX1 \FIFO_reg[50][24]  ( .D(n2955), .CLK(clk_in), .RSTB(n7195), .Q(
        \FIFO[50][24] ) );
  DFFARX1 \FIFO_reg[50][23]  ( .D(n2954), .CLK(clk_in), .RSTB(n7196), .Q(
        \FIFO[50][23] ) );
  DFFARX1 \FIFO_reg[50][22]  ( .D(n2953), .CLK(clk_in), .RSTB(n7196), .Q(
        \FIFO[50][22] ) );
  DFFARX1 \FIFO_reg[50][21]  ( .D(n2952), .CLK(clk_in), .RSTB(n7196), .Q(
        \FIFO[50][21] ) );
  DFFARX1 \FIFO_reg[50][20]  ( .D(n2951), .CLK(clk_in), .RSTB(n7196), .Q(
        \FIFO[50][20] ) );
  DFFARX1 \FIFO_reg[50][19]  ( .D(n2950), .CLK(clk_in), .RSTB(n7196), .Q(
        \FIFO[50][19] ) );
  DFFARX1 \FIFO_reg[50][18]  ( .D(n2949), .CLK(clk_in), .RSTB(n7196), .Q(
        \FIFO[50][18] ) );
  DFFARX1 \FIFO_reg[50][17]  ( .D(n2948), .CLK(clk_in), .RSTB(n7196), .Q(
        \FIFO[50][17] ) );
  DFFARX1 \FIFO_reg[50][16]  ( .D(n2947), .CLK(clk_in), .RSTB(n7196), .Q(
        \FIFO[50][16] ) );
  DFFARX1 \FIFO_reg[50][15]  ( .D(n2946), .CLK(clk_in), .RSTB(n7196), .Q(
        \FIFO[50][15] ) );
  DFFARX1 \FIFO_reg[50][14]  ( .D(n2945), .CLK(clk_in), .RSTB(n7196), .Q(
        \FIFO[50][14] ) );
  DFFARX1 \FIFO_reg[50][13]  ( .D(n2944), .CLK(clk_in), .RSTB(n7196), .Q(
        \FIFO[50][13] ) );
  DFFARX1 \FIFO_reg[50][12]  ( .D(n2943), .CLK(clk_in), .RSTB(n7196), .Q(
        \FIFO[50][12] ) );
  DFFARX1 \FIFO_reg[50][11]  ( .D(n2942), .CLK(clk_in), .RSTB(n7196), .Q(
        \FIFO[50][11] ) );
  DFFARX1 \FIFO_reg[50][10]  ( .D(n2941), .CLK(clk_in), .RSTB(n7196), .Q(
        \FIFO[50][10] ) );
  DFFARX1 \FIFO_reg[50][9]  ( .D(n2940), .CLK(clk_in), .RSTB(n7196), .Q(
        \FIFO[50][9] ) );
  DFFARX1 \FIFO_reg[50][8]  ( .D(n2939), .CLK(clk_in), .RSTB(n7196), .Q(
        \FIFO[50][8] ) );
  DFFARX1 \FIFO_reg[50][7]  ( .D(n2938), .CLK(clk_in), .RSTB(n7196), .Q(
        \FIFO[50][7] ) );
  DFFARX1 \FIFO_reg[50][6]  ( .D(n2937), .CLK(clk_in), .RSTB(n7196), .Q(
        \FIFO[50][6] ) );
  DFFARX1 \FIFO_reg[50][5]  ( .D(n2936), .CLK(clk_in), .RSTB(n7197), .Q(
        \FIFO[50][5] ) );
  DFFARX1 \FIFO_reg[50][4]  ( .D(n2935), .CLK(clk_in), .RSTB(n7197), .Q(
        \FIFO[50][4] ) );
  DFFARX1 \FIFO_reg[50][3]  ( .D(n2934), .CLK(clk_in), .RSTB(n7197), .Q(
        \FIFO[50][3] ) );
  DFFARX1 \FIFO_reg[50][2]  ( .D(n2933), .CLK(clk_in), .RSTB(n7197), .Q(
        \FIFO[50][2] ) );
  DFFARX1 \FIFO_reg[50][1]  ( .D(n2932), .CLK(clk_in), .RSTB(n7197), .Q(
        \FIFO[50][1] ) );
  DFFARX1 \FIFO_reg[50][0]  ( .D(n2931), .CLK(clk_in), .RSTB(n7197), .Q(
        \FIFO[50][0] ) );
  DFFARX1 \FIFO_reg[51][31]  ( .D(n2930), .CLK(clk_in), .RSTB(n7197), .Q(
        \FIFO[51][31] ) );
  DFFARX1 \FIFO_reg[51][30]  ( .D(n2929), .CLK(clk_in), .RSTB(n7197), .Q(
        \FIFO[51][30] ) );
  DFFARX1 \FIFO_reg[51][29]  ( .D(n2928), .CLK(clk_in), .RSTB(n7197), .Q(
        \FIFO[51][29] ) );
  DFFARX1 \FIFO_reg[51][28]  ( .D(n2927), .CLK(clk_in), .RSTB(n7197), .Q(
        \FIFO[51][28] ) );
  DFFARX1 \FIFO_reg[51][27]  ( .D(n2926), .CLK(clk_in), .RSTB(n7197), .Q(
        \FIFO[51][27] ) );
  DFFARX1 \FIFO_reg[51][26]  ( .D(n2925), .CLK(clk_in), .RSTB(n7197), .Q(
        \FIFO[51][26] ) );
  DFFARX1 \FIFO_reg[51][25]  ( .D(n2924), .CLK(clk_in), .RSTB(n7197), .Q(
        \FIFO[51][25] ) );
  DFFARX1 \FIFO_reg[51][24]  ( .D(n2923), .CLK(clk_in), .RSTB(n7197), .Q(
        \FIFO[51][24] ) );
  DFFARX1 \FIFO_reg[51][23]  ( .D(n2922), .CLK(clk_in), .RSTB(n7197), .Q(
        \FIFO[51][23] ) );
  DFFARX1 \FIFO_reg[51][22]  ( .D(n2921), .CLK(clk_in), .RSTB(n7197), .Q(
        \FIFO[51][22] ) );
  DFFARX1 \FIFO_reg[51][21]  ( .D(n2920), .CLK(clk_in), .RSTB(n7197), .Q(
        \FIFO[51][21] ) );
  DFFARX1 \FIFO_reg[51][20]  ( .D(n2919), .CLK(clk_in), .RSTB(n7197), .Q(
        \FIFO[51][20] ) );
  DFFARX1 \FIFO_reg[51][19]  ( .D(n2918), .CLK(clk_in), .RSTB(n7198), .Q(
        \FIFO[51][19] ) );
  DFFARX1 \FIFO_reg[51][18]  ( .D(n2917), .CLK(clk_in), .RSTB(n7198), .Q(
        \FIFO[51][18] ) );
  DFFARX1 \FIFO_reg[51][17]  ( .D(n2916), .CLK(clk_in), .RSTB(n7198), .Q(
        \FIFO[51][17] ) );
  DFFARX1 \FIFO_reg[51][16]  ( .D(n2915), .CLK(clk_in), .RSTB(n7198), .Q(
        \FIFO[51][16] ) );
  DFFARX1 \FIFO_reg[51][15]  ( .D(n2914), .CLK(clk_in), .RSTB(n7198), .Q(
        \FIFO[51][15] ) );
  DFFARX1 \FIFO_reg[51][14]  ( .D(n2913), .CLK(clk_in), .RSTB(n7198), .Q(
        \FIFO[51][14] ) );
  DFFARX1 \FIFO_reg[51][13]  ( .D(n2912), .CLK(clk_in), .RSTB(n7198), .Q(
        \FIFO[51][13] ) );
  DFFARX1 \FIFO_reg[51][12]  ( .D(n2911), .CLK(clk_in), .RSTB(n7198), .Q(
        \FIFO[51][12] ) );
  DFFARX1 \FIFO_reg[51][11]  ( .D(n2910), .CLK(clk_in), .RSTB(n7198), .Q(
        \FIFO[51][11] ) );
  DFFARX1 \FIFO_reg[51][10]  ( .D(n2909), .CLK(clk_in), .RSTB(n7198), .Q(
        \FIFO[51][10] ) );
  DFFARX1 \FIFO_reg[51][9]  ( .D(n2908), .CLK(clk_in), .RSTB(n7198), .Q(
        \FIFO[51][9] ) );
  DFFARX1 \FIFO_reg[51][8]  ( .D(n2907), .CLK(clk_in), .RSTB(n7198), .Q(
        \FIFO[51][8] ) );
  DFFARX1 \FIFO_reg[51][7]  ( .D(n2906), .CLK(clk_in), .RSTB(n7198), .Q(
        \FIFO[51][7] ) );
  DFFARX1 \FIFO_reg[51][6]  ( .D(n2905), .CLK(clk_in), .RSTB(n7198), .Q(
        \FIFO[51][6] ) );
  DFFARX1 \FIFO_reg[51][5]  ( .D(n2904), .CLK(clk_in), .RSTB(n7198), .Q(
        \FIFO[51][5] ) );
  DFFARX1 \FIFO_reg[51][4]  ( .D(n2903), .CLK(clk_in), .RSTB(n7198), .Q(
        \FIFO[51][4] ) );
  DFFARX1 \FIFO_reg[51][3]  ( .D(n2902), .CLK(clk_in), .RSTB(n7198), .Q(
        \FIFO[51][3] ) );
  DFFARX1 \FIFO_reg[51][2]  ( .D(n2901), .CLK(clk_in), .RSTB(n7198), .Q(
        \FIFO[51][2] ) );
  DFFARX1 \FIFO_reg[51][1]  ( .D(n2900), .CLK(clk_in), .RSTB(n7199), .Q(
        \FIFO[51][1] ) );
  DFFARX1 \FIFO_reg[51][0]  ( .D(n2899), .CLK(clk_in), .RSTB(n7199), .Q(
        \FIFO[51][0] ) );
  DFFARX1 \FIFO_reg[52][31]  ( .D(n2898), .CLK(clk_in), .RSTB(n7199), .Q(
        \FIFO[52][31] ) );
  DFFARX1 \FIFO_reg[52][30]  ( .D(n2897), .CLK(clk_in), .RSTB(n7199), .Q(
        \FIFO[52][30] ) );
  DFFARX1 \FIFO_reg[52][29]  ( .D(n2896), .CLK(clk_in), .RSTB(n7199), .Q(
        \FIFO[52][29] ) );
  DFFARX1 \FIFO_reg[52][28]  ( .D(n2895), .CLK(clk_in), .RSTB(n7199), .Q(
        \FIFO[52][28] ) );
  DFFARX1 \FIFO_reg[52][27]  ( .D(n2894), .CLK(clk_in), .RSTB(n7199), .Q(
        \FIFO[52][27] ) );
  DFFARX1 \FIFO_reg[52][26]  ( .D(n2893), .CLK(clk_in), .RSTB(n7199), .Q(
        \FIFO[52][26] ) );
  DFFARX1 \FIFO_reg[52][25]  ( .D(n2892), .CLK(clk_in), .RSTB(n7199), .Q(
        \FIFO[52][25] ) );
  DFFARX1 \FIFO_reg[52][24]  ( .D(n2891), .CLK(clk_in), .RSTB(n7199), .Q(
        \FIFO[52][24] ) );
  DFFARX1 \FIFO_reg[52][23]  ( .D(n2890), .CLK(clk_in), .RSTB(n7199), .Q(
        \FIFO[52][23] ) );
  DFFARX1 \FIFO_reg[52][22]  ( .D(n2889), .CLK(clk_in), .RSTB(n7199), .Q(
        \FIFO[52][22] ) );
  DFFARX1 \FIFO_reg[52][21]  ( .D(n2888), .CLK(clk_in), .RSTB(n7199), .Q(
        \FIFO[52][21] ) );
  DFFARX1 \FIFO_reg[52][20]  ( .D(n2887), .CLK(clk_in), .RSTB(n7199), .Q(
        \FIFO[52][20] ) );
  DFFARX1 \FIFO_reg[52][19]  ( .D(n2886), .CLK(clk_in), .RSTB(n7199), .Q(
        \FIFO[52][19] ) );
  DFFARX1 \FIFO_reg[52][18]  ( .D(n2885), .CLK(clk_in), .RSTB(n7199), .Q(
        \FIFO[52][18] ) );
  DFFARX1 \FIFO_reg[52][17]  ( .D(n2884), .CLK(clk_in), .RSTB(n7199), .Q(
        \FIFO[52][17] ) );
  DFFARX1 \FIFO_reg[52][16]  ( .D(n2883), .CLK(clk_in), .RSTB(n7199), .Q(
        \FIFO[52][16] ) );
  DFFARX1 \FIFO_reg[52][15]  ( .D(n2882), .CLK(clk_in), .RSTB(n7200), .Q(
        \FIFO[52][15] ) );
  DFFARX1 \FIFO_reg[52][14]  ( .D(n2881), .CLK(clk_in), .RSTB(n7200), .Q(
        \FIFO[52][14] ) );
  DFFARX1 \FIFO_reg[52][13]  ( .D(n2880), .CLK(clk_in), .RSTB(n7200), .Q(
        \FIFO[52][13] ) );
  DFFARX1 \FIFO_reg[52][12]  ( .D(n2879), .CLK(clk_in), .RSTB(n7200), .Q(
        \FIFO[52][12] ) );
  DFFARX1 \FIFO_reg[52][11]  ( .D(n2878), .CLK(clk_in), .RSTB(n7200), .Q(
        \FIFO[52][11] ) );
  DFFARX1 \FIFO_reg[52][10]  ( .D(n2877), .CLK(clk_in), .RSTB(n7200), .Q(
        \FIFO[52][10] ) );
  DFFARX1 \FIFO_reg[52][9]  ( .D(n2876), .CLK(clk_in), .RSTB(n7200), .Q(
        \FIFO[52][9] ) );
  DFFARX1 \FIFO_reg[52][8]  ( .D(n2875), .CLK(clk_in), .RSTB(n7200), .Q(
        \FIFO[52][8] ) );
  DFFARX1 \FIFO_reg[52][7]  ( .D(n2874), .CLK(clk_in), .RSTB(n7200), .Q(
        \FIFO[52][7] ) );
  DFFARX1 \FIFO_reg[52][6]  ( .D(n2873), .CLK(clk_in), .RSTB(n7200), .Q(
        \FIFO[52][6] ) );
  DFFARX1 \FIFO_reg[52][5]  ( .D(n2872), .CLK(clk_in), .RSTB(n7200), .Q(
        \FIFO[52][5] ) );
  DFFARX1 \FIFO_reg[52][4]  ( .D(n2871), .CLK(clk_in), .RSTB(n7200), .Q(
        \FIFO[52][4] ) );
  DFFARX1 \FIFO_reg[52][3]  ( .D(n2870), .CLK(clk_in), .RSTB(n7200), .Q(
        \FIFO[52][3] ) );
  DFFARX1 \FIFO_reg[52][2]  ( .D(n2869), .CLK(clk_in), .RSTB(n7200), .Q(
        \FIFO[52][2] ) );
  DFFARX1 \FIFO_reg[52][1]  ( .D(n2868), .CLK(clk_in), .RSTB(n7200), .Q(
        \FIFO[52][1] ) );
  DFFARX1 \FIFO_reg[52][0]  ( .D(n2867), .CLK(clk_in), .RSTB(n7200), .Q(
        \FIFO[52][0] ) );
  DFFARX1 \FIFO_reg[53][31]  ( .D(n2866), .CLK(clk_in), .RSTB(n7200), .Q(
        \FIFO[53][31] ) );
  DFFARX1 \FIFO_reg[53][30]  ( .D(n2865), .CLK(clk_in), .RSTB(n7200), .Q(
        \FIFO[53][30] ) );
  DFFARX1 \FIFO_reg[53][29]  ( .D(n2864), .CLK(clk_in), .RSTB(n7201), .Q(
        \FIFO[53][29] ) );
  DFFARX1 \FIFO_reg[53][28]  ( .D(n2863), .CLK(clk_in), .RSTB(n7201), .Q(
        \FIFO[53][28] ) );
  DFFARX1 \FIFO_reg[53][27]  ( .D(n2862), .CLK(clk_in), .RSTB(n7201), .Q(
        \FIFO[53][27] ) );
  DFFARX1 \FIFO_reg[53][26]  ( .D(n2861), .CLK(clk_in), .RSTB(n7201), .Q(
        \FIFO[53][26] ) );
  DFFARX1 \FIFO_reg[53][25]  ( .D(n2860), .CLK(clk_in), .RSTB(n7201), .Q(
        \FIFO[53][25] ) );
  DFFARX1 \FIFO_reg[53][24]  ( .D(n2859), .CLK(clk_in), .RSTB(n7201), .Q(
        \FIFO[53][24] ) );
  DFFARX1 \FIFO_reg[53][23]  ( .D(n2858), .CLK(clk_in), .RSTB(n7201), .Q(
        \FIFO[53][23] ) );
  DFFARX1 \FIFO_reg[53][22]  ( .D(n2857), .CLK(clk_in), .RSTB(n7201), .Q(
        \FIFO[53][22] ) );
  DFFARX1 \FIFO_reg[53][21]  ( .D(n2856), .CLK(clk_in), .RSTB(n7201), .Q(
        \FIFO[53][21] ) );
  DFFARX1 \FIFO_reg[53][20]  ( .D(n2855), .CLK(clk_in), .RSTB(n7201), .Q(
        \FIFO[53][20] ) );
  DFFARX1 \FIFO_reg[53][19]  ( .D(n2854), .CLK(clk_in), .RSTB(n7201), .Q(
        \FIFO[53][19] ) );
  DFFARX1 \FIFO_reg[53][18]  ( .D(n2853), .CLK(clk_in), .RSTB(n7201), .Q(
        \FIFO[53][18] ) );
  DFFARX1 \FIFO_reg[53][17]  ( .D(n2852), .CLK(clk_in), .RSTB(n7201), .Q(
        \FIFO[53][17] ) );
  DFFARX1 \FIFO_reg[53][16]  ( .D(n2851), .CLK(clk_in), .RSTB(n7201), .Q(
        \FIFO[53][16] ) );
  DFFARX1 \FIFO_reg[53][15]  ( .D(n2850), .CLK(clk_in), .RSTB(n7201), .Q(
        \FIFO[53][15] ) );
  DFFARX1 \FIFO_reg[53][14]  ( .D(n2849), .CLK(clk_in), .RSTB(n7201), .Q(
        \FIFO[53][14] ) );
  DFFARX1 \FIFO_reg[53][13]  ( .D(n2848), .CLK(clk_in), .RSTB(n7201), .Q(
        \FIFO[53][13] ) );
  DFFARX1 \FIFO_reg[53][12]  ( .D(n2847), .CLK(clk_in), .RSTB(n7201), .Q(
        \FIFO[53][12] ) );
  DFFARX1 \FIFO_reg[53][11]  ( .D(n2846), .CLK(clk_in), .RSTB(n7202), .Q(
        \FIFO[53][11] ) );
  DFFARX1 \FIFO_reg[53][10]  ( .D(n2845), .CLK(clk_in), .RSTB(n7202), .Q(
        \FIFO[53][10] ) );
  DFFARX1 \FIFO_reg[53][9]  ( .D(n2844), .CLK(clk_in), .RSTB(n7202), .Q(
        \FIFO[53][9] ) );
  DFFARX1 \FIFO_reg[53][8]  ( .D(n2843), .CLK(clk_in), .RSTB(n7202), .Q(
        \FIFO[53][8] ) );
  DFFARX1 \FIFO_reg[53][7]  ( .D(n2842), .CLK(clk_in), .RSTB(n7202), .Q(
        \FIFO[53][7] ) );
  DFFARX1 \FIFO_reg[53][6]  ( .D(n2841), .CLK(clk_in), .RSTB(n7202), .Q(
        \FIFO[53][6] ) );
  DFFARX1 \FIFO_reg[53][5]  ( .D(n2840), .CLK(clk_in), .RSTB(n7202), .Q(
        \FIFO[53][5] ) );
  DFFARX1 \FIFO_reg[53][4]  ( .D(n2839), .CLK(clk_in), .RSTB(n7202), .Q(
        \FIFO[53][4] ) );
  DFFARX1 \FIFO_reg[53][3]  ( .D(n2838), .CLK(clk_in), .RSTB(n7202), .Q(
        \FIFO[53][3] ) );
  DFFARX1 \FIFO_reg[53][2]  ( .D(n2837), .CLK(clk_in), .RSTB(n7202), .Q(
        \FIFO[53][2] ) );
  DFFARX1 \FIFO_reg[53][1]  ( .D(n2836), .CLK(clk_in), .RSTB(n7202), .Q(
        \FIFO[53][1] ) );
  DFFARX1 \FIFO_reg[53][0]  ( .D(n2835), .CLK(clk_in), .RSTB(n7202), .Q(
        \FIFO[53][0] ) );
  DFFARX1 \FIFO_reg[54][31]  ( .D(n2834), .CLK(clk_in), .RSTB(n7202), .Q(
        \FIFO[54][31] ) );
  DFFARX1 \FIFO_reg[54][30]  ( .D(n2833), .CLK(clk_in), .RSTB(n7202), .Q(
        \FIFO[54][30] ) );
  DFFARX1 \FIFO_reg[54][29]  ( .D(n2832), .CLK(clk_in), .RSTB(n7202), .Q(
        \FIFO[54][29] ) );
  DFFARX1 \FIFO_reg[54][28]  ( .D(n2831), .CLK(clk_in), .RSTB(n7202), .Q(
        \FIFO[54][28] ) );
  DFFARX1 \FIFO_reg[54][27]  ( .D(n2830), .CLK(clk_in), .RSTB(n7202), .Q(
        \FIFO[54][27] ) );
  DFFARX1 \FIFO_reg[54][26]  ( .D(n2829), .CLK(clk_in), .RSTB(n7202), .Q(
        \FIFO[54][26] ) );
  DFFARX1 \FIFO_reg[54][25]  ( .D(n2828), .CLK(clk_in), .RSTB(n7203), .Q(
        \FIFO[54][25] ) );
  DFFARX1 \FIFO_reg[54][24]  ( .D(n2827), .CLK(clk_in), .RSTB(n7203), .Q(
        \FIFO[54][24] ) );
  DFFARX1 \FIFO_reg[54][23]  ( .D(n2826), .CLK(clk_in), .RSTB(n7203), .Q(
        \FIFO[54][23] ) );
  DFFARX1 \FIFO_reg[54][22]  ( .D(n2825), .CLK(clk_in), .RSTB(n7203), .Q(
        \FIFO[54][22] ) );
  DFFARX1 \FIFO_reg[54][21]  ( .D(n2824), .CLK(clk_in), .RSTB(n7203), .Q(
        \FIFO[54][21] ) );
  DFFARX1 \FIFO_reg[54][20]  ( .D(n2823), .CLK(clk_in), .RSTB(n7203), .Q(
        \FIFO[54][20] ) );
  DFFARX1 \FIFO_reg[54][19]  ( .D(n2822), .CLK(clk_in), .RSTB(n7203), .Q(
        \FIFO[54][19] ) );
  DFFARX1 \FIFO_reg[54][18]  ( .D(n2821), .CLK(clk_in), .RSTB(n7203), .Q(
        \FIFO[54][18] ) );
  DFFARX1 \FIFO_reg[54][17]  ( .D(n2820), .CLK(clk_in), .RSTB(n7203), .Q(
        \FIFO[54][17] ) );
  DFFARX1 \FIFO_reg[54][16]  ( .D(n2819), .CLK(clk_in), .RSTB(n7203), .Q(
        \FIFO[54][16] ) );
  DFFARX1 \FIFO_reg[54][15]  ( .D(n2818), .CLK(clk_in), .RSTB(n7203), .Q(
        \FIFO[54][15] ) );
  DFFARX1 \FIFO_reg[54][14]  ( .D(n2817), .CLK(clk_in), .RSTB(n7203), .Q(
        \FIFO[54][14] ) );
  DFFARX1 \FIFO_reg[54][13]  ( .D(n2816), .CLK(clk_in), .RSTB(n7203), .Q(
        \FIFO[54][13] ) );
  DFFARX1 \FIFO_reg[54][12]  ( .D(n2815), .CLK(clk_in), .RSTB(n7203), .Q(
        \FIFO[54][12] ) );
  DFFARX1 \FIFO_reg[54][11]  ( .D(n2814), .CLK(clk_in), .RSTB(n7203), .Q(
        \FIFO[54][11] ) );
  DFFARX1 \FIFO_reg[54][10]  ( .D(n2813), .CLK(clk_in), .RSTB(n7203), .Q(
        \FIFO[54][10] ) );
  DFFARX1 \FIFO_reg[54][9]  ( .D(n2812), .CLK(clk_in), .RSTB(n7203), .Q(
        \FIFO[54][9] ) );
  DFFARX1 \FIFO_reg[54][8]  ( .D(n2811), .CLK(clk_in), .RSTB(n7203), .Q(
        \FIFO[54][8] ) );
  DFFARX1 \FIFO_reg[54][7]  ( .D(n2810), .CLK(clk_in), .RSTB(n7204), .Q(
        \FIFO[54][7] ) );
  DFFARX1 \FIFO_reg[54][6]  ( .D(n2809), .CLK(clk_in), .RSTB(n7204), .Q(
        \FIFO[54][6] ) );
  DFFARX1 \FIFO_reg[54][5]  ( .D(n2808), .CLK(clk_in), .RSTB(n7204), .Q(
        \FIFO[54][5] ) );
  DFFARX1 \FIFO_reg[54][4]  ( .D(n2807), .CLK(clk_in), .RSTB(n7204), .Q(
        \FIFO[54][4] ) );
  DFFARX1 \FIFO_reg[54][3]  ( .D(n2806), .CLK(clk_in), .RSTB(n7204), .Q(
        \FIFO[54][3] ) );
  DFFARX1 \FIFO_reg[54][2]  ( .D(n2805), .CLK(clk_in), .RSTB(n7204), .Q(
        \FIFO[54][2] ) );
  DFFARX1 \FIFO_reg[54][1]  ( .D(n2804), .CLK(clk_in), .RSTB(n7204), .Q(
        \FIFO[54][1] ) );
  DFFARX1 \FIFO_reg[54][0]  ( .D(n2803), .CLK(clk_in), .RSTB(n7204), .Q(
        \FIFO[54][0] ) );
  DFFARX1 \FIFO_reg[55][31]  ( .D(n2802), .CLK(clk_in), .RSTB(n7204), .Q(
        \FIFO[55][31] ) );
  DFFARX1 \FIFO_reg[55][30]  ( .D(n2801), .CLK(clk_in), .RSTB(n7204), .Q(
        \FIFO[55][30] ) );
  DFFARX1 \FIFO_reg[55][29]  ( .D(n2800), .CLK(clk_in), .RSTB(n7204), .Q(
        \FIFO[55][29] ) );
  DFFARX1 \FIFO_reg[55][28]  ( .D(n2799), .CLK(clk_in), .RSTB(n7204), .Q(
        \FIFO[55][28] ) );
  DFFARX1 \FIFO_reg[55][27]  ( .D(n2798), .CLK(clk_in), .RSTB(n7204), .Q(
        \FIFO[55][27] ) );
  DFFARX1 \FIFO_reg[55][26]  ( .D(n2797), .CLK(clk_in), .RSTB(n7204), .Q(
        \FIFO[55][26] ) );
  DFFARX1 \FIFO_reg[55][25]  ( .D(n2796), .CLK(clk_in), .RSTB(n7204), .Q(
        \FIFO[55][25] ) );
  DFFARX1 \FIFO_reg[55][24]  ( .D(n2795), .CLK(clk_in), .RSTB(n7204), .Q(
        \FIFO[55][24] ) );
  DFFARX1 \FIFO_reg[55][23]  ( .D(n2794), .CLK(clk_in), .RSTB(n7204), .Q(
        \FIFO[55][23] ) );
  DFFARX1 \FIFO_reg[55][22]  ( .D(n2793), .CLK(clk_in), .RSTB(n7204), .Q(
        \FIFO[55][22] ) );
  DFFARX1 \FIFO_reg[55][21]  ( .D(n2792), .CLK(clk_in), .RSTB(n7205), .Q(
        \FIFO[55][21] ) );
  DFFARX1 \FIFO_reg[55][20]  ( .D(n2791), .CLK(clk_in), .RSTB(n7205), .Q(
        \FIFO[55][20] ) );
  DFFARX1 \FIFO_reg[55][19]  ( .D(n2790), .CLK(clk_in), .RSTB(n7205), .Q(
        \FIFO[55][19] ) );
  DFFARX1 \FIFO_reg[55][18]  ( .D(n2789), .CLK(clk_in), .RSTB(n7205), .Q(
        \FIFO[55][18] ) );
  DFFARX1 \FIFO_reg[55][17]  ( .D(n2788), .CLK(clk_in), .RSTB(n7205), .Q(
        \FIFO[55][17] ) );
  DFFARX1 \FIFO_reg[55][16]  ( .D(n2787), .CLK(clk_in), .RSTB(n7205), .Q(
        \FIFO[55][16] ) );
  DFFARX1 \FIFO_reg[55][15]  ( .D(n2786), .CLK(clk_in), .RSTB(n7205), .Q(
        \FIFO[55][15] ) );
  DFFARX1 \FIFO_reg[55][14]  ( .D(n2785), .CLK(clk_in), .RSTB(n7205), .Q(
        \FIFO[55][14] ) );
  DFFARX1 \FIFO_reg[55][13]  ( .D(n2784), .CLK(clk_in), .RSTB(n7205), .Q(
        \FIFO[55][13] ) );
  DFFARX1 \FIFO_reg[55][12]  ( .D(n2783), .CLK(clk_in), .RSTB(n7205), .Q(
        \FIFO[55][12] ) );
  DFFARX1 \FIFO_reg[55][11]  ( .D(n2782), .CLK(clk_in), .RSTB(n7205), .Q(
        \FIFO[55][11] ) );
  DFFARX1 \FIFO_reg[55][10]  ( .D(n2781), .CLK(clk_in), .RSTB(n7205), .Q(
        \FIFO[55][10] ) );
  DFFARX1 \FIFO_reg[55][9]  ( .D(n2780), .CLK(clk_in), .RSTB(n7205), .Q(
        \FIFO[55][9] ) );
  DFFARX1 \FIFO_reg[55][8]  ( .D(n2779), .CLK(clk_in), .RSTB(n7205), .Q(
        \FIFO[55][8] ) );
  DFFARX1 \FIFO_reg[55][7]  ( .D(n2778), .CLK(clk_in), .RSTB(n7205), .Q(
        \FIFO[55][7] ) );
  DFFARX1 \FIFO_reg[55][6]  ( .D(n2777), .CLK(clk_in), .RSTB(n7205), .Q(
        \FIFO[55][6] ) );
  DFFARX1 \FIFO_reg[55][5]  ( .D(n2776), .CLK(clk_in), .RSTB(n7205), .Q(
        \FIFO[55][5] ) );
  DFFARX1 \FIFO_reg[55][4]  ( .D(n2775), .CLK(clk_in), .RSTB(n7205), .Q(
        \FIFO[55][4] ) );
  DFFARX1 \FIFO_reg[55][3]  ( .D(n2774), .CLK(clk_in), .RSTB(n7206), .Q(
        \FIFO[55][3] ) );
  DFFARX1 \FIFO_reg[55][2]  ( .D(n2773), .CLK(clk_in), .RSTB(n7206), .Q(
        \FIFO[55][2] ) );
  DFFARX1 \FIFO_reg[55][1]  ( .D(n2772), .CLK(clk_in), .RSTB(n7206), .Q(
        \FIFO[55][1] ) );
  DFFARX1 \FIFO_reg[55][0]  ( .D(n2771), .CLK(clk_in), .RSTB(n7206), .Q(
        \FIFO[55][0] ) );
  DFFARX1 \FIFO_reg[56][31]  ( .D(n2770), .CLK(clk_in), .RSTB(n7206), .Q(
        \FIFO[56][31] ) );
  DFFARX1 \FIFO_reg[56][30]  ( .D(n2769), .CLK(clk_in), .RSTB(n7206), .Q(
        \FIFO[56][30] ) );
  DFFARX1 \FIFO_reg[56][29]  ( .D(n2768), .CLK(clk_in), .RSTB(n7206), .Q(
        \FIFO[56][29] ) );
  DFFARX1 \FIFO_reg[56][28]  ( .D(n2767), .CLK(clk_in), .RSTB(n7206), .Q(
        \FIFO[56][28] ) );
  DFFARX1 \FIFO_reg[56][27]  ( .D(n2766), .CLK(clk_in), .RSTB(n7206), .Q(
        \FIFO[56][27] ) );
  DFFARX1 \FIFO_reg[56][26]  ( .D(n2765), .CLK(clk_in), .RSTB(n7206), .Q(
        \FIFO[56][26] ) );
  DFFARX1 \FIFO_reg[56][25]  ( .D(n2764), .CLK(clk_in), .RSTB(n7206), .Q(
        \FIFO[56][25] ) );
  DFFARX1 \FIFO_reg[56][24]  ( .D(n2763), .CLK(clk_in), .RSTB(n7206), .Q(
        \FIFO[56][24] ) );
  DFFARX1 \FIFO_reg[56][23]  ( .D(n2762), .CLK(clk_in), .RSTB(n7206), .Q(
        \FIFO[56][23] ) );
  DFFARX1 \FIFO_reg[56][22]  ( .D(n2761), .CLK(clk_in), .RSTB(n7206), .Q(
        \FIFO[56][22] ) );
  DFFARX1 \FIFO_reg[56][21]  ( .D(n2760), .CLK(clk_in), .RSTB(n7206), .Q(
        \FIFO[56][21] ) );
  DFFARX1 \FIFO_reg[56][20]  ( .D(n2759), .CLK(clk_in), .RSTB(n7206), .Q(
        \FIFO[56][20] ) );
  DFFARX1 \FIFO_reg[56][19]  ( .D(n2758), .CLK(clk_in), .RSTB(n7206), .Q(
        \FIFO[56][19] ) );
  DFFARX1 \FIFO_reg[56][18]  ( .D(n2757), .CLK(clk_in), .RSTB(n7206), .Q(
        \FIFO[56][18] ) );
  DFFARX1 \FIFO_reg[56][17]  ( .D(n2756), .CLK(clk_in), .RSTB(n7207), .Q(
        \FIFO[56][17] ) );
  DFFARX1 \FIFO_reg[56][16]  ( .D(n2755), .CLK(clk_in), .RSTB(n7207), .Q(
        \FIFO[56][16] ) );
  DFFARX1 \FIFO_reg[56][15]  ( .D(n2754), .CLK(clk_in), .RSTB(n7207), .Q(
        \FIFO[56][15] ) );
  DFFARX1 \FIFO_reg[56][14]  ( .D(n2753), .CLK(clk_in), .RSTB(n7207), .Q(
        \FIFO[56][14] ) );
  DFFARX1 \FIFO_reg[56][13]  ( .D(n2752), .CLK(clk_in), .RSTB(n7207), .Q(
        \FIFO[56][13] ) );
  DFFARX1 \FIFO_reg[56][12]  ( .D(n2751), .CLK(clk_in), .RSTB(n7207), .Q(
        \FIFO[56][12] ) );
  DFFARX1 \FIFO_reg[56][11]  ( .D(n2750), .CLK(clk_in), .RSTB(n7207), .Q(
        \FIFO[56][11] ) );
  DFFARX1 \FIFO_reg[56][10]  ( .D(n2749), .CLK(clk_in), .RSTB(n7207), .Q(
        \FIFO[56][10] ) );
  DFFARX1 \FIFO_reg[56][9]  ( .D(n2748), .CLK(clk_in), .RSTB(n7207), .Q(
        \FIFO[56][9] ) );
  DFFARX1 \FIFO_reg[56][8]  ( .D(n2747), .CLK(clk_in), .RSTB(n7207), .Q(
        \FIFO[56][8] ) );
  DFFARX1 \FIFO_reg[56][7]  ( .D(n2746), .CLK(clk_in), .RSTB(n7207), .Q(
        \FIFO[56][7] ) );
  DFFARX1 \FIFO_reg[56][6]  ( .D(n2745), .CLK(clk_in), .RSTB(n7207), .Q(
        \FIFO[56][6] ) );
  DFFARX1 \FIFO_reg[56][5]  ( .D(n2744), .CLK(clk_in), .RSTB(n7207), .Q(
        \FIFO[56][5] ) );
  DFFARX1 \FIFO_reg[56][4]  ( .D(n2743), .CLK(clk_in), .RSTB(n7207), .Q(
        \FIFO[56][4] ) );
  DFFARX1 \FIFO_reg[56][3]  ( .D(n2742), .CLK(clk_in), .RSTB(n7207), .Q(
        \FIFO[56][3] ) );
  DFFARX1 \FIFO_reg[56][2]  ( .D(n2741), .CLK(clk_in), .RSTB(n7207), .Q(
        \FIFO[56][2] ) );
  DFFARX1 \FIFO_reg[56][1]  ( .D(n2740), .CLK(clk_in), .RSTB(n7207), .Q(
        \FIFO[56][1] ) );
  DFFARX1 \FIFO_reg[56][0]  ( .D(n2739), .CLK(clk_in), .RSTB(n7207), .Q(
        \FIFO[56][0] ) );
  DFFARX1 \FIFO_reg[57][31]  ( .D(n2738), .CLK(clk_in), .RSTB(n7208), .Q(
        \FIFO[57][31] ) );
  DFFARX1 \FIFO_reg[57][30]  ( .D(n2737), .CLK(clk_in), .RSTB(n7208), .Q(
        \FIFO[57][30] ) );
  DFFARX1 \FIFO_reg[57][29]  ( .D(n2736), .CLK(clk_in), .RSTB(n7208), .Q(
        \FIFO[57][29] ) );
  DFFARX1 \FIFO_reg[57][28]  ( .D(n2735), .CLK(clk_in), .RSTB(n7208), .Q(
        \FIFO[57][28] ) );
  DFFARX1 \FIFO_reg[57][27]  ( .D(n2734), .CLK(clk_in), .RSTB(n7208), .Q(
        \FIFO[57][27] ) );
  DFFARX1 \FIFO_reg[57][26]  ( .D(n2733), .CLK(clk_in), .RSTB(n7208), .Q(
        \FIFO[57][26] ) );
  DFFARX1 \FIFO_reg[57][25]  ( .D(n2732), .CLK(clk_in), .RSTB(n7208), .Q(
        \FIFO[57][25] ) );
  DFFARX1 \FIFO_reg[57][24]  ( .D(n2731), .CLK(clk_in), .RSTB(n7208), .Q(
        \FIFO[57][24] ) );
  DFFARX1 \FIFO_reg[57][23]  ( .D(n2730), .CLK(clk_in), .RSTB(n7208), .Q(
        \FIFO[57][23] ) );
  DFFARX1 \FIFO_reg[57][22]  ( .D(n2729), .CLK(clk_in), .RSTB(n7208), .Q(
        \FIFO[57][22] ) );
  DFFARX1 \FIFO_reg[57][21]  ( .D(n2728), .CLK(clk_in), .RSTB(n7208), .Q(
        \FIFO[57][21] ) );
  DFFARX1 \FIFO_reg[57][20]  ( .D(n2727), .CLK(clk_in), .RSTB(n7208), .Q(
        \FIFO[57][20] ) );
  DFFARX1 \FIFO_reg[57][19]  ( .D(n2726), .CLK(clk_in), .RSTB(n7208), .Q(
        \FIFO[57][19] ) );
  DFFARX1 \FIFO_reg[57][18]  ( .D(n2725), .CLK(clk_in), .RSTB(n7208), .Q(
        \FIFO[57][18] ) );
  DFFARX1 \FIFO_reg[57][17]  ( .D(n2724), .CLK(clk_in), .RSTB(n7208), .Q(
        \FIFO[57][17] ) );
  DFFARX1 \FIFO_reg[57][16]  ( .D(n2723), .CLK(clk_in), .RSTB(n7208), .Q(
        \FIFO[57][16] ) );
  DFFARX1 \FIFO_reg[57][15]  ( .D(n2722), .CLK(clk_in), .RSTB(n7208), .Q(
        \FIFO[57][15] ) );
  DFFARX1 \FIFO_reg[57][14]  ( .D(n2721), .CLK(clk_in), .RSTB(n7208), .Q(
        \FIFO[57][14] ) );
  DFFARX1 \FIFO_reg[57][13]  ( .D(n2720), .CLK(clk_in), .RSTB(n7209), .Q(
        \FIFO[57][13] ) );
  DFFARX1 \FIFO_reg[57][12]  ( .D(n2719), .CLK(clk_in), .RSTB(n7209), .Q(
        \FIFO[57][12] ) );
  DFFARX1 \FIFO_reg[57][11]  ( .D(n2718), .CLK(clk_in), .RSTB(n7209), .Q(
        \FIFO[57][11] ) );
  DFFARX1 \FIFO_reg[57][10]  ( .D(n2717), .CLK(clk_in), .RSTB(n7209), .Q(
        \FIFO[57][10] ) );
  DFFARX1 \FIFO_reg[57][9]  ( .D(n2716), .CLK(clk_in), .RSTB(n7209), .Q(
        \FIFO[57][9] ) );
  DFFARX1 \FIFO_reg[57][8]  ( .D(n2715), .CLK(clk_in), .RSTB(n7209), .Q(
        \FIFO[57][8] ) );
  DFFARX1 \FIFO_reg[57][7]  ( .D(n2714), .CLK(clk_in), .RSTB(n7209), .Q(
        \FIFO[57][7] ) );
  DFFARX1 \FIFO_reg[57][6]  ( .D(n2713), .CLK(clk_in), .RSTB(n7209), .Q(
        \FIFO[57][6] ) );
  DFFARX1 \FIFO_reg[57][5]  ( .D(n2712), .CLK(clk_in), .RSTB(n7209), .Q(
        \FIFO[57][5] ) );
  DFFARX1 \FIFO_reg[57][4]  ( .D(n2711), .CLK(clk_in), .RSTB(n7209), .Q(
        \FIFO[57][4] ) );
  DFFARX1 \FIFO_reg[57][3]  ( .D(n2710), .CLK(clk_in), .RSTB(n7209), .Q(
        \FIFO[57][3] ) );
  DFFARX1 \FIFO_reg[57][2]  ( .D(n2709), .CLK(clk_in), .RSTB(n7209), .Q(
        \FIFO[57][2] ) );
  DFFARX1 \FIFO_reg[57][1]  ( .D(n2708), .CLK(clk_in), .RSTB(n7209), .Q(
        \FIFO[57][1] ) );
  DFFARX1 \FIFO_reg[57][0]  ( .D(n2707), .CLK(clk_in), .RSTB(n7209), .Q(
        \FIFO[57][0] ) );
  DFFARX1 \FIFO_reg[58][31]  ( .D(n2706), .CLK(clk_in), .RSTB(n7209), .Q(
        \FIFO[58][31] ) );
  DFFARX1 \FIFO_reg[58][30]  ( .D(n2705), .CLK(clk_in), .RSTB(n7209), .Q(
        \FIFO[58][30] ) );
  DFFARX1 \FIFO_reg[58][29]  ( .D(n2704), .CLK(clk_in), .RSTB(n7209), .Q(
        \FIFO[58][29] ) );
  DFFARX1 \FIFO_reg[58][28]  ( .D(n2703), .CLK(clk_in), .RSTB(n7209), .Q(
        \FIFO[58][28] ) );
  DFFARX1 \FIFO_reg[58][27]  ( .D(n2702), .CLK(clk_in), .RSTB(n7210), .Q(
        \FIFO[58][27] ) );
  DFFARX1 \FIFO_reg[58][26]  ( .D(n2701), .CLK(clk_in), .RSTB(n7210), .Q(
        \FIFO[58][26] ) );
  DFFARX1 \FIFO_reg[58][25]  ( .D(n2700), .CLK(clk_in), .RSTB(n7210), .Q(
        \FIFO[58][25] ) );
  DFFARX1 \FIFO_reg[58][24]  ( .D(n2699), .CLK(clk_in), .RSTB(n7210), .Q(
        \FIFO[58][24] ) );
  DFFARX1 \FIFO_reg[58][23]  ( .D(n2698), .CLK(clk_in), .RSTB(n7210), .Q(
        \FIFO[58][23] ) );
  DFFARX1 \FIFO_reg[58][22]  ( .D(n2697), .CLK(clk_in), .RSTB(n7210), .Q(
        \FIFO[58][22] ) );
  DFFARX1 \FIFO_reg[58][21]  ( .D(n2696), .CLK(clk_in), .RSTB(n7210), .Q(
        \FIFO[58][21] ) );
  DFFARX1 \FIFO_reg[58][20]  ( .D(n2695), .CLK(clk_in), .RSTB(n7210), .Q(
        \FIFO[58][20] ) );
  DFFARX1 \FIFO_reg[58][19]  ( .D(n2694), .CLK(clk_in), .RSTB(n7210), .Q(
        \FIFO[58][19] ) );
  DFFARX1 \FIFO_reg[58][18]  ( .D(n2693), .CLK(clk_in), .RSTB(n7210), .Q(
        \FIFO[58][18] ) );
  DFFARX1 \FIFO_reg[58][17]  ( .D(n2692), .CLK(clk_in), .RSTB(n7210), .Q(
        \FIFO[58][17] ) );
  DFFARX1 \FIFO_reg[58][16]  ( .D(n2691), .CLK(clk_in), .RSTB(n7210), .Q(
        \FIFO[58][16] ) );
  DFFARX1 \FIFO_reg[58][15]  ( .D(n2690), .CLK(clk_in), .RSTB(n7210), .Q(
        \FIFO[58][15] ) );
  DFFARX1 \FIFO_reg[58][14]  ( .D(n2689), .CLK(clk_in), .RSTB(n7210), .Q(
        \FIFO[58][14] ) );
  DFFARX1 \FIFO_reg[58][13]  ( .D(n2688), .CLK(clk_in), .RSTB(n7210), .Q(
        \FIFO[58][13] ) );
  DFFARX1 \FIFO_reg[58][12]  ( .D(n2687), .CLK(clk_in), .RSTB(n7210), .Q(
        \FIFO[58][12] ) );
  DFFARX1 \FIFO_reg[58][11]  ( .D(n2686), .CLK(clk_in), .RSTB(n7210), .Q(
        \FIFO[58][11] ) );
  DFFARX1 \FIFO_reg[58][10]  ( .D(n2685), .CLK(clk_in), .RSTB(n7210), .Q(
        \FIFO[58][10] ) );
  DFFARX1 \FIFO_reg[58][9]  ( .D(n2684), .CLK(clk_in), .RSTB(n7211), .Q(
        \FIFO[58][9] ) );
  DFFARX1 \FIFO_reg[58][8]  ( .D(n2683), .CLK(clk_in), .RSTB(n7211), .Q(
        \FIFO[58][8] ) );
  DFFARX1 \FIFO_reg[58][7]  ( .D(n2682), .CLK(clk_in), .RSTB(n7211), .Q(
        \FIFO[58][7] ) );
  DFFARX1 \FIFO_reg[58][6]  ( .D(n2681), .CLK(clk_in), .RSTB(n7211), .Q(
        \FIFO[58][6] ) );
  DFFARX1 \FIFO_reg[58][5]  ( .D(n2680), .CLK(clk_in), .RSTB(n7211), .Q(
        \FIFO[58][5] ) );
  DFFARX1 \FIFO_reg[58][4]  ( .D(n2679), .CLK(clk_in), .RSTB(n7211), .Q(
        \FIFO[58][4] ) );
  DFFARX1 \FIFO_reg[58][3]  ( .D(n2678), .CLK(clk_in), .RSTB(n7211), .Q(
        \FIFO[58][3] ) );
  DFFARX1 \FIFO_reg[58][2]  ( .D(n2677), .CLK(clk_in), .RSTB(n7211), .Q(
        \FIFO[58][2] ) );
  DFFARX1 \FIFO_reg[58][1]  ( .D(n2676), .CLK(clk_in), .RSTB(n7211), .Q(
        \FIFO[58][1] ) );
  DFFARX1 \FIFO_reg[58][0]  ( .D(n2675), .CLK(clk_in), .RSTB(n7211), .Q(
        \FIFO[58][0] ) );
  DFFARX1 \FIFO_reg[59][31]  ( .D(n2674), .CLK(clk_in), .RSTB(n7211), .Q(
        \FIFO[59][31] ) );
  DFFARX1 \FIFO_reg[59][30]  ( .D(n2673), .CLK(clk_in), .RSTB(n7211), .Q(
        \FIFO[59][30] ) );
  DFFARX1 \FIFO_reg[59][29]  ( .D(n2672), .CLK(clk_in), .RSTB(n7211), .Q(
        \FIFO[59][29] ) );
  DFFARX1 \FIFO_reg[59][28]  ( .D(n2671), .CLK(clk_in), .RSTB(n7211), .Q(
        \FIFO[59][28] ) );
  DFFARX1 \FIFO_reg[59][27]  ( .D(n2670), .CLK(clk_in), .RSTB(n7211), .Q(
        \FIFO[59][27] ) );
  DFFARX1 \FIFO_reg[59][26]  ( .D(n2669), .CLK(clk_in), .RSTB(n7211), .Q(
        \FIFO[59][26] ) );
  DFFARX1 \FIFO_reg[59][25]  ( .D(n2668), .CLK(clk_in), .RSTB(n7211), .Q(
        \FIFO[59][25] ) );
  DFFARX1 \FIFO_reg[59][24]  ( .D(n2667), .CLK(clk_in), .RSTB(n7211), .Q(
        \FIFO[59][24] ) );
  DFFARX1 \FIFO_reg[59][23]  ( .D(n2666), .CLK(clk_in), .RSTB(n7212), .Q(
        \FIFO[59][23] ) );
  DFFARX1 \FIFO_reg[59][22]  ( .D(n2665), .CLK(clk_in), .RSTB(n7212), .Q(
        \FIFO[59][22] ) );
  DFFARX1 \FIFO_reg[59][21]  ( .D(n2664), .CLK(clk_in), .RSTB(n7212), .Q(
        \FIFO[59][21] ) );
  DFFARX1 \FIFO_reg[59][20]  ( .D(n2663), .CLK(clk_in), .RSTB(n7212), .Q(
        \FIFO[59][20] ) );
  DFFARX1 \FIFO_reg[59][19]  ( .D(n2662), .CLK(clk_in), .RSTB(n7212), .Q(
        \FIFO[59][19] ) );
  DFFARX1 \FIFO_reg[59][18]  ( .D(n2661), .CLK(clk_in), .RSTB(n7212), .Q(
        \FIFO[59][18] ) );
  DFFARX1 \FIFO_reg[59][17]  ( .D(n2660), .CLK(clk_in), .RSTB(n7212), .Q(
        \FIFO[59][17] ) );
  DFFARX1 \FIFO_reg[59][16]  ( .D(n2659), .CLK(clk_in), .RSTB(n7212), .Q(
        \FIFO[59][16] ) );
  DFFARX1 \FIFO_reg[59][15]  ( .D(n2658), .CLK(clk_in), .RSTB(n7212), .Q(
        \FIFO[59][15] ) );
  DFFARX1 \FIFO_reg[59][14]  ( .D(n2657), .CLK(clk_in), .RSTB(n7212), .Q(
        \FIFO[59][14] ) );
  DFFARX1 \FIFO_reg[59][13]  ( .D(n2656), .CLK(clk_in), .RSTB(n7212), .Q(
        \FIFO[59][13] ) );
  DFFARX1 \FIFO_reg[59][12]  ( .D(n2655), .CLK(clk_in), .RSTB(n7212), .Q(
        \FIFO[59][12] ) );
  DFFARX1 \FIFO_reg[59][11]  ( .D(n2654), .CLK(clk_in), .RSTB(n7212), .Q(
        \FIFO[59][11] ) );
  DFFARX1 \FIFO_reg[59][10]  ( .D(n2653), .CLK(clk_in), .RSTB(n7212), .Q(
        \FIFO[59][10] ) );
  DFFARX1 \FIFO_reg[59][9]  ( .D(n2652), .CLK(clk_in), .RSTB(n7212), .Q(
        \FIFO[59][9] ) );
  DFFARX1 \FIFO_reg[59][8]  ( .D(n2651), .CLK(clk_in), .RSTB(n7212), .Q(
        \FIFO[59][8] ) );
  DFFARX1 \FIFO_reg[59][7]  ( .D(n2650), .CLK(clk_in), .RSTB(n7212), .Q(
        \FIFO[59][7] ) );
  DFFARX1 \FIFO_reg[59][6]  ( .D(n2649), .CLK(clk_in), .RSTB(n7212), .Q(
        \FIFO[59][6] ) );
  DFFARX1 \FIFO_reg[59][5]  ( .D(n2648), .CLK(clk_in), .RSTB(n7213), .Q(
        \FIFO[59][5] ) );
  DFFARX1 \FIFO_reg[59][4]  ( .D(n2647), .CLK(clk_in), .RSTB(n7213), .Q(
        \FIFO[59][4] ) );
  DFFARX1 \FIFO_reg[59][3]  ( .D(n2646), .CLK(clk_in), .RSTB(n7213), .Q(
        \FIFO[59][3] ) );
  DFFARX1 \FIFO_reg[59][2]  ( .D(n2645), .CLK(clk_in), .RSTB(n7213), .Q(
        \FIFO[59][2] ) );
  DFFARX1 \FIFO_reg[59][1]  ( .D(n2644), .CLK(clk_in), .RSTB(n7213), .Q(
        \FIFO[59][1] ) );
  DFFARX1 \FIFO_reg[59][0]  ( .D(n2643), .CLK(clk_in), .RSTB(n7213), .Q(
        \FIFO[59][0] ) );
  DFFARX1 \FIFO_reg[60][31]  ( .D(n2642), .CLK(clk_in), .RSTB(n7213), .Q(
        \FIFO[60][31] ) );
  DFFARX1 \FIFO_reg[60][30]  ( .D(n2641), .CLK(clk_in), .RSTB(n7213), .Q(
        \FIFO[60][30] ) );
  DFFARX1 \FIFO_reg[60][29]  ( .D(n2640), .CLK(clk_in), .RSTB(n7213), .Q(
        \FIFO[60][29] ) );
  DFFARX1 \FIFO_reg[60][28]  ( .D(n2639), .CLK(clk_in), .RSTB(n7213), .Q(
        \FIFO[60][28] ) );
  DFFARX1 \FIFO_reg[60][27]  ( .D(n2638), .CLK(clk_in), .RSTB(n7213), .Q(
        \FIFO[60][27] ) );
  DFFARX1 \FIFO_reg[60][26]  ( .D(n2637), .CLK(clk_in), .RSTB(n7213), .Q(
        \FIFO[60][26] ) );
  DFFARX1 \FIFO_reg[60][25]  ( .D(n2636), .CLK(clk_in), .RSTB(n7213), .Q(
        \FIFO[60][25] ) );
  DFFARX1 \FIFO_reg[60][24]  ( .D(n2635), .CLK(clk_in), .RSTB(n7213), .Q(
        \FIFO[60][24] ) );
  DFFARX1 \FIFO_reg[60][23]  ( .D(n2634), .CLK(clk_in), .RSTB(n7213), .Q(
        \FIFO[60][23] ) );
  DFFARX1 \FIFO_reg[60][22]  ( .D(n2633), .CLK(clk_in), .RSTB(n7213), .Q(
        \FIFO[60][22] ) );
  DFFARX1 \FIFO_reg[60][21]  ( .D(n2632), .CLK(clk_in), .RSTB(n7213), .Q(
        \FIFO[60][21] ) );
  DFFARX1 \FIFO_reg[60][20]  ( .D(n2631), .CLK(clk_in), .RSTB(n7213), .Q(
        \FIFO[60][20] ) );
  DFFARX1 \FIFO_reg[60][19]  ( .D(n2630), .CLK(clk_in), .RSTB(n7214), .Q(
        \FIFO[60][19] ) );
  DFFARX1 \FIFO_reg[60][18]  ( .D(n2629), .CLK(clk_in), .RSTB(n7214), .Q(
        \FIFO[60][18] ) );
  DFFARX1 \FIFO_reg[60][17]  ( .D(n2628), .CLK(clk_in), .RSTB(n7214), .Q(
        \FIFO[60][17] ) );
  DFFARX1 \FIFO_reg[60][16]  ( .D(n2627), .CLK(clk_in), .RSTB(n7214), .Q(
        \FIFO[60][16] ) );
  DFFARX1 \FIFO_reg[60][15]  ( .D(n2626), .CLK(clk_in), .RSTB(n7214), .Q(
        \FIFO[60][15] ) );
  DFFARX1 \FIFO_reg[60][14]  ( .D(n2625), .CLK(clk_in), .RSTB(n7214), .Q(
        \FIFO[60][14] ) );
  DFFARX1 \FIFO_reg[60][13]  ( .D(n2624), .CLK(clk_in), .RSTB(n7214), .Q(
        \FIFO[60][13] ) );
  DFFARX1 \FIFO_reg[60][12]  ( .D(n2623), .CLK(clk_in), .RSTB(n7214), .Q(
        \FIFO[60][12] ) );
  DFFARX1 \FIFO_reg[60][11]  ( .D(n2622), .CLK(clk_in), .RSTB(n7214), .Q(
        \FIFO[60][11] ) );
  DFFARX1 \FIFO_reg[60][10]  ( .D(n2621), .CLK(clk_in), .RSTB(n7214), .Q(
        \FIFO[60][10] ) );
  DFFARX1 \FIFO_reg[60][9]  ( .D(n2620), .CLK(clk_in), .RSTB(n7214), .Q(
        \FIFO[60][9] ) );
  DFFARX1 \FIFO_reg[60][8]  ( .D(n2619), .CLK(clk_in), .RSTB(n7214), .Q(
        \FIFO[60][8] ) );
  DFFARX1 \FIFO_reg[60][7]  ( .D(n2618), .CLK(clk_in), .RSTB(n7214), .Q(
        \FIFO[60][7] ) );
  DFFARX1 \FIFO_reg[60][6]  ( .D(n2617), .CLK(clk_in), .RSTB(n7214), .Q(
        \FIFO[60][6] ) );
  DFFARX1 \FIFO_reg[60][5]  ( .D(n2616), .CLK(clk_in), .RSTB(n7214), .Q(
        \FIFO[60][5] ) );
  DFFARX1 \FIFO_reg[60][4]  ( .D(n2615), .CLK(clk_in), .RSTB(n7214), .Q(
        \FIFO[60][4] ) );
  DFFARX1 \FIFO_reg[60][3]  ( .D(n2614), .CLK(clk_in), .RSTB(n7214), .Q(
        \FIFO[60][3] ) );
  DFFARX1 \FIFO_reg[60][2]  ( .D(n2613), .CLK(clk_in), .RSTB(n7214), .Q(
        \FIFO[60][2] ) );
  DFFARX1 \FIFO_reg[60][1]  ( .D(n2612), .CLK(clk_in), .RSTB(n7215), .Q(
        \FIFO[60][1] ) );
  DFFARX1 \FIFO_reg[60][0]  ( .D(n2611), .CLK(clk_in), .RSTB(n7215), .Q(
        \FIFO[60][0] ) );
  DFFARX1 \FIFO_reg[61][31]  ( .D(n2610), .CLK(clk_in), .RSTB(n7215), .Q(
        \FIFO[61][31] ) );
  DFFARX1 \FIFO_reg[61][30]  ( .D(n2609), .CLK(clk_in), .RSTB(n7215), .Q(
        \FIFO[61][30] ) );
  DFFARX1 \FIFO_reg[61][29]  ( .D(n2608), .CLK(clk_in), .RSTB(n7215), .Q(
        \FIFO[61][29] ) );
  DFFARX1 \FIFO_reg[61][28]  ( .D(n2607), .CLK(clk_in), .RSTB(n7215), .Q(
        \FIFO[61][28] ) );
  DFFARX1 \FIFO_reg[61][27]  ( .D(n2606), .CLK(clk_in), .RSTB(n7215), .Q(
        \FIFO[61][27] ) );
  DFFARX1 \FIFO_reg[61][26]  ( .D(n2605), .CLK(clk_in), .RSTB(n7215), .Q(
        \FIFO[61][26] ) );
  DFFARX1 \FIFO_reg[61][25]  ( .D(n2604), .CLK(clk_in), .RSTB(n7215), .Q(
        \FIFO[61][25] ) );
  DFFARX1 \FIFO_reg[61][24]  ( .D(n2603), .CLK(clk_in), .RSTB(n7215), .Q(
        \FIFO[61][24] ) );
  DFFARX1 \FIFO_reg[61][23]  ( .D(n2602), .CLK(clk_in), .RSTB(n7215), .Q(
        \FIFO[61][23] ) );
  DFFARX1 \FIFO_reg[61][22]  ( .D(n2601), .CLK(clk_in), .RSTB(n7215), .Q(
        \FIFO[61][22] ) );
  DFFARX1 \FIFO_reg[61][21]  ( .D(n2600), .CLK(clk_in), .RSTB(n7215), .Q(
        \FIFO[61][21] ) );
  DFFARX1 \FIFO_reg[61][20]  ( .D(n2599), .CLK(clk_in), .RSTB(n7215), .Q(
        \FIFO[61][20] ) );
  DFFARX1 \FIFO_reg[61][19]  ( .D(n2598), .CLK(clk_in), .RSTB(n7215), .Q(
        \FIFO[61][19] ) );
  DFFARX1 \FIFO_reg[61][18]  ( .D(n2597), .CLK(clk_in), .RSTB(n7215), .Q(
        \FIFO[61][18] ) );
  DFFARX1 \FIFO_reg[61][17]  ( .D(n2596), .CLK(clk_in), .RSTB(n7215), .Q(
        \FIFO[61][17] ) );
  DFFARX1 \FIFO_reg[61][16]  ( .D(n2595), .CLK(clk_in), .RSTB(n7215), .Q(
        \FIFO[61][16] ) );
  DFFARX1 \FIFO_reg[61][15]  ( .D(n2594), .CLK(clk_in), .RSTB(n7216), .Q(
        \FIFO[61][15] ) );
  DFFARX1 \FIFO_reg[61][14]  ( .D(n2593), .CLK(clk_in), .RSTB(n7216), .Q(
        \FIFO[61][14] ) );
  DFFARX1 \FIFO_reg[61][13]  ( .D(n2592), .CLK(clk_in), .RSTB(n7216), .Q(
        \FIFO[61][13] ) );
  DFFARX1 \FIFO_reg[61][12]  ( .D(n2591), .CLK(clk_in), .RSTB(n7216), .Q(
        \FIFO[61][12] ) );
  DFFARX1 \FIFO_reg[61][11]  ( .D(n2590), .CLK(clk_in), .RSTB(n7216), .Q(
        \FIFO[61][11] ) );
  DFFARX1 \FIFO_reg[61][10]  ( .D(n2589), .CLK(clk_in), .RSTB(n7216), .Q(
        \FIFO[61][10] ) );
  DFFARX1 \FIFO_reg[61][9]  ( .D(n2588), .CLK(clk_in), .RSTB(n7216), .Q(
        \FIFO[61][9] ) );
  DFFARX1 \FIFO_reg[61][8]  ( .D(n2587), .CLK(clk_in), .RSTB(n7216), .Q(
        \FIFO[61][8] ) );
  DFFARX1 \FIFO_reg[61][7]  ( .D(n2586), .CLK(clk_in), .RSTB(n7216), .Q(
        \FIFO[61][7] ) );
  DFFARX1 \FIFO_reg[61][6]  ( .D(n2585), .CLK(clk_in), .RSTB(n7216), .Q(
        \FIFO[61][6] ) );
  DFFARX1 \FIFO_reg[61][5]  ( .D(n2584), .CLK(clk_in), .RSTB(n7216), .Q(
        \FIFO[61][5] ) );
  DFFARX1 \FIFO_reg[61][4]  ( .D(n2583), .CLK(clk_in), .RSTB(n7216), .Q(
        \FIFO[61][4] ) );
  DFFARX1 \FIFO_reg[61][3]  ( .D(n2582), .CLK(clk_in), .RSTB(n7216), .Q(
        \FIFO[61][3] ) );
  DFFARX1 \FIFO_reg[61][2]  ( .D(n2581), .CLK(clk_in), .RSTB(n7216), .Q(
        \FIFO[61][2] ) );
  DFFARX1 \FIFO_reg[61][1]  ( .D(n2580), .CLK(clk_in), .RSTB(n7216), .Q(
        \FIFO[61][1] ) );
  DFFARX1 \FIFO_reg[61][0]  ( .D(n2579), .CLK(clk_in), .RSTB(n7216), .Q(
        \FIFO[61][0] ) );
  DFFARX1 \FIFO_reg[62][31]  ( .D(n2578), .CLK(clk_in), .RSTB(n7216), .Q(
        \FIFO[62][31] ) );
  DFFARX1 \FIFO_reg[62][30]  ( .D(n2577), .CLK(clk_in), .RSTB(n7216), .Q(
        \FIFO[62][30] ) );
  DFFARX1 \FIFO_reg[62][29]  ( .D(n2576), .CLK(clk_in), .RSTB(n7217), .Q(
        \FIFO[62][29] ) );
  DFFARX1 \FIFO_reg[62][28]  ( .D(n2575), .CLK(clk_in), .RSTB(n7217), .Q(
        \FIFO[62][28] ) );
  DFFARX1 \FIFO_reg[62][27]  ( .D(n2574), .CLK(clk_in), .RSTB(n7217), .Q(
        \FIFO[62][27] ) );
  DFFARX1 \FIFO_reg[62][26]  ( .D(n2573), .CLK(clk_in), .RSTB(n7217), .Q(
        \FIFO[62][26] ) );
  DFFARX1 \FIFO_reg[62][25]  ( .D(n2572), .CLK(clk_in), .RSTB(n7217), .Q(
        \FIFO[62][25] ) );
  DFFARX1 \FIFO_reg[62][24]  ( .D(n2571), .CLK(clk_in), .RSTB(n7217), .Q(
        \FIFO[62][24] ) );
  DFFARX1 \FIFO_reg[62][23]  ( .D(n2570), .CLK(clk_in), .RSTB(n7217), .Q(
        \FIFO[62][23] ) );
  DFFARX1 \FIFO_reg[62][22]  ( .D(n2569), .CLK(clk_in), .RSTB(n7217), .Q(
        \FIFO[62][22] ) );
  DFFARX1 \FIFO_reg[62][21]  ( .D(n2568), .CLK(clk_in), .RSTB(n7217), .Q(
        \FIFO[62][21] ) );
  DFFARX1 \FIFO_reg[62][20]  ( .D(n2567), .CLK(clk_in), .RSTB(n7217), .Q(
        \FIFO[62][20] ) );
  DFFARX1 \FIFO_reg[62][19]  ( .D(n2566), .CLK(clk_in), .RSTB(n7217), .Q(
        \FIFO[62][19] ) );
  DFFARX1 \FIFO_reg[62][18]  ( .D(n2565), .CLK(clk_in), .RSTB(n7217), .Q(
        \FIFO[62][18] ) );
  DFFARX1 \FIFO_reg[62][17]  ( .D(n2564), .CLK(clk_in), .RSTB(n7217), .Q(
        \FIFO[62][17] ) );
  DFFARX1 \FIFO_reg[62][16]  ( .D(n2563), .CLK(clk_in), .RSTB(n7217), .Q(
        \FIFO[62][16] ) );
  DFFARX1 \FIFO_reg[62][15]  ( .D(n2562), .CLK(clk_in), .RSTB(n7217), .Q(
        \FIFO[62][15] ) );
  DFFARX1 \FIFO_reg[62][14]  ( .D(n2561), .CLK(clk_in), .RSTB(n7217), .Q(
        \FIFO[62][14] ) );
  DFFARX1 \FIFO_reg[62][13]  ( .D(n2560), .CLK(clk_in), .RSTB(n7217), .Q(
        \FIFO[62][13] ) );
  DFFARX1 \FIFO_reg[62][12]  ( .D(n2559), .CLK(clk_in), .RSTB(n7217), .Q(
        \FIFO[62][12] ) );
  DFFARX1 \FIFO_reg[62][11]  ( .D(n2558), .CLK(clk_in), .RSTB(n7218), .Q(
        \FIFO[62][11] ) );
  DFFARX1 \FIFO_reg[62][10]  ( .D(n2557), .CLK(clk_in), .RSTB(n7218), .Q(
        \FIFO[62][10] ) );
  DFFARX1 \FIFO_reg[62][9]  ( .D(n2556), .CLK(clk_in), .RSTB(n7218), .Q(
        \FIFO[62][9] ) );
  DFFARX1 \FIFO_reg[62][8]  ( .D(n2555), .CLK(clk_in), .RSTB(n7218), .Q(
        \FIFO[62][8] ) );
  DFFARX1 \FIFO_reg[62][7]  ( .D(n2554), .CLK(clk_in), .RSTB(n7218), .Q(
        \FIFO[62][7] ) );
  DFFARX1 \FIFO_reg[62][6]  ( .D(n2553), .CLK(clk_in), .RSTB(n7218), .Q(
        \FIFO[62][6] ) );
  DFFARX1 \FIFO_reg[62][5]  ( .D(n2552), .CLK(clk_in), .RSTB(n7218), .Q(
        \FIFO[62][5] ) );
  DFFARX1 \FIFO_reg[62][4]  ( .D(n2551), .CLK(clk_in), .RSTB(n7218), .Q(
        \FIFO[62][4] ) );
  DFFARX1 \FIFO_reg[62][3]  ( .D(n2550), .CLK(clk_in), .RSTB(n7218), .Q(
        \FIFO[62][3] ) );
  DFFARX1 \FIFO_reg[62][2]  ( .D(n2549), .CLK(clk_in), .RSTB(n7218), .Q(
        \FIFO[62][2] ) );
  DFFARX1 \FIFO_reg[62][1]  ( .D(n2548), .CLK(clk_in), .RSTB(n7218), .Q(
        \FIFO[62][1] ) );
  DFFARX1 \FIFO_reg[62][0]  ( .D(n2547), .CLK(clk_in), .RSTB(n7218), .Q(
        \FIFO[62][0] ) );
  DFFARX1 \FIFO_reg[63][31]  ( .D(n2546), .CLK(clk_in), .RSTB(n7218), .Q(
        \FIFO[63][31] ) );
  DFFARX1 \FIFO_reg[63][30]  ( .D(n2545), .CLK(clk_in), .RSTB(n7218), .Q(
        \FIFO[63][30] ) );
  DFFARX1 \FIFO_reg[63][29]  ( .D(n2544), .CLK(clk_in), .RSTB(n7218), .Q(
        \FIFO[63][29] ) );
  DFFARX1 \FIFO_reg[63][28]  ( .D(n2543), .CLK(clk_in), .RSTB(n7218), .Q(
        \FIFO[63][28] ) );
  DFFARX1 \FIFO_reg[63][27]  ( .D(n2542), .CLK(clk_in), .RSTB(n7218), .Q(
        \FIFO[63][27] ) );
  DFFARX1 \FIFO_reg[63][26]  ( .D(n2541), .CLK(clk_in), .RSTB(n7218), .Q(
        \FIFO[63][26] ) );
  DFFARX1 \FIFO_reg[63][25]  ( .D(n2540), .CLK(clk_in), .RSTB(n7219), .Q(
        \FIFO[63][25] ) );
  DFFARX1 \FIFO_reg[63][24]  ( .D(n2539), .CLK(clk_in), .RSTB(n7219), .Q(
        \FIFO[63][24] ) );
  DFFARX1 \FIFO_reg[63][23]  ( .D(n2538), .CLK(clk_in), .RSTB(n7219), .Q(
        \FIFO[63][23] ) );
  DFFARX1 \FIFO_reg[63][22]  ( .D(n2537), .CLK(clk_in), .RSTB(n7219), .Q(
        \FIFO[63][22] ) );
  DFFARX1 \FIFO_reg[63][21]  ( .D(n2536), .CLK(clk_in), .RSTB(n7219), .Q(
        \FIFO[63][21] ) );
  DFFARX1 \FIFO_reg[63][20]  ( .D(n2535), .CLK(clk_in), .RSTB(n7219), .Q(
        \FIFO[63][20] ) );
  DFFARX1 \FIFO_reg[63][19]  ( .D(n2534), .CLK(clk_in), .RSTB(n7219), .Q(
        \FIFO[63][19] ) );
  DFFARX1 \FIFO_reg[63][18]  ( .D(n2533), .CLK(clk_in), .RSTB(n7219), .Q(
        \FIFO[63][18] ) );
  DFFARX1 \FIFO_reg[63][17]  ( .D(n2532), .CLK(clk_in), .RSTB(n7219), .Q(
        \FIFO[63][17] ) );
  DFFARX1 \FIFO_reg[63][16]  ( .D(n2531), .CLK(clk_in), .RSTB(n7219), .Q(
        \FIFO[63][16] ) );
  DFFARX1 \FIFO_reg[63][15]  ( .D(n2530), .CLK(clk_in), .RSTB(n7219), .Q(
        \FIFO[63][15] ) );
  DFFARX1 \FIFO_reg[63][14]  ( .D(n2529), .CLK(clk_in), .RSTB(n7219), .Q(
        \FIFO[63][14] ) );
  DFFARX1 \FIFO_reg[63][13]  ( .D(n2528), .CLK(clk_in), .RSTB(n7219), .Q(
        \FIFO[63][13] ) );
  DFFARX1 \FIFO_reg[63][12]  ( .D(n2527), .CLK(clk_in), .RSTB(n7219), .Q(
        \FIFO[63][12] ) );
  DFFARX1 \FIFO_reg[63][11]  ( .D(n2526), .CLK(clk_in), .RSTB(n7219), .Q(
        \FIFO[63][11] ) );
  DFFARX1 \FIFO_reg[63][10]  ( .D(n2525), .CLK(clk_in), .RSTB(n7219), .Q(
        \FIFO[63][10] ) );
  DFFARX1 \FIFO_reg[63][9]  ( .D(n2524), .CLK(clk_in), .RSTB(n7219), .Q(
        \FIFO[63][9] ) );
  DFFARX1 \FIFO_reg[63][8]  ( .D(n2523), .CLK(clk_in), .RSTB(n7219), .Q(
        \FIFO[63][8] ) );
  DFFARX1 \FIFO_reg[63][7]  ( .D(n2522), .CLK(clk_in), .RSTB(n7220), .Q(
        \FIFO[63][7] ) );
  DFFARX1 \FIFO_reg[63][6]  ( .D(n2521), .CLK(clk_in), .RSTB(n7220), .Q(
        \FIFO[63][6] ) );
  DFFARX1 \FIFO_reg[63][5]  ( .D(n2520), .CLK(clk_in), .RSTB(n7220), .Q(
        \FIFO[63][5] ) );
  DFFARX1 \FIFO_reg[63][4]  ( .D(n2519), .CLK(clk_in), .RSTB(n7220), .Q(
        \FIFO[63][4] ) );
  DFFARX1 \FIFO_reg[63][3]  ( .D(n2518), .CLK(clk_in), .RSTB(n7220), .Q(
        \FIFO[63][3] ) );
  DFFARX1 \FIFO_reg[63][2]  ( .D(n2517), .CLK(clk_in), .RSTB(n7220), .Q(
        \FIFO[63][2] ) );
  DFFARX1 \FIFO_reg[63][1]  ( .D(n2516), .CLK(clk_in), .RSTB(n7220), .Q(
        \FIFO[63][1] ) );
  DFFARX1 \FIFO_reg[63][0]  ( .D(n2515), .CLK(clk_in), .RSTB(n7220), .Q(
        \FIFO[63][0] ) );
  DFFARX1 \FIFO_reg[64][31]  ( .D(n2514), .CLK(clk_in), .RSTB(n7220), .Q(
        \FIFO[64][31] ) );
  DFFARX1 \FIFO_reg[64][30]  ( .D(n2513), .CLK(clk_in), .RSTB(n7220), .Q(
        \FIFO[64][30] ) );
  DFFARX1 \FIFO_reg[64][29]  ( .D(n2512), .CLK(clk_in), .RSTB(n7220), .Q(
        \FIFO[64][29] ) );
  DFFARX1 \FIFO_reg[64][28]  ( .D(n2511), .CLK(clk_in), .RSTB(n7220), .Q(
        \FIFO[64][28] ) );
  DFFARX1 \FIFO_reg[64][27]  ( .D(n2510), .CLK(clk_in), .RSTB(n7220), .Q(
        \FIFO[64][27] ) );
  DFFARX1 \FIFO_reg[64][26]  ( .D(n2509), .CLK(clk_in), .RSTB(n7220), .Q(
        \FIFO[64][26] ) );
  DFFARX1 \FIFO_reg[64][25]  ( .D(n2508), .CLK(clk_in), .RSTB(n7220), .Q(
        \FIFO[64][25] ) );
  DFFARX1 \FIFO_reg[64][24]  ( .D(n2507), .CLK(clk_in), .RSTB(n7220), .Q(
        \FIFO[64][24] ) );
  DFFARX1 \FIFO_reg[64][23]  ( .D(n2506), .CLK(clk_in), .RSTB(n7220), .Q(
        \FIFO[64][23] ) );
  DFFARX1 \FIFO_reg[64][22]  ( .D(n2505), .CLK(clk_in), .RSTB(n7220), .Q(
        \FIFO[64][22] ) );
  DFFARX1 \FIFO_reg[64][21]  ( .D(n2504), .CLK(clk_in), .RSTB(n7221), .Q(
        \FIFO[64][21] ) );
  DFFARX1 \FIFO_reg[64][20]  ( .D(n2503), .CLK(clk_in), .RSTB(n7221), .Q(
        \FIFO[64][20] ) );
  DFFARX1 \FIFO_reg[64][19]  ( .D(n2502), .CLK(clk_in), .RSTB(n7221), .Q(
        \FIFO[64][19] ) );
  DFFARX1 \FIFO_reg[64][18]  ( .D(n2501), .CLK(clk_in), .RSTB(n7221), .Q(
        \FIFO[64][18] ) );
  DFFARX1 \FIFO_reg[64][17]  ( .D(n2500), .CLK(clk_in), .RSTB(n7221), .Q(
        \FIFO[64][17] ) );
  DFFARX1 \FIFO_reg[64][16]  ( .D(n2499), .CLK(clk_in), .RSTB(n7221), .Q(
        \FIFO[64][16] ) );
  DFFARX1 \FIFO_reg[64][15]  ( .D(n2498), .CLK(clk_in), .RSTB(n7221), .Q(
        \FIFO[64][15] ) );
  DFFARX1 \FIFO_reg[64][14]  ( .D(n2497), .CLK(clk_in), .RSTB(n7221), .Q(
        \FIFO[64][14] ) );
  DFFARX1 \FIFO_reg[64][13]  ( .D(n2496), .CLK(clk_in), .RSTB(n7221), .Q(
        \FIFO[64][13] ) );
  DFFARX1 \FIFO_reg[64][12]  ( .D(n2495), .CLK(clk_in), .RSTB(n7221), .Q(
        \FIFO[64][12] ) );
  DFFARX1 \FIFO_reg[64][11]  ( .D(n2494), .CLK(clk_in), .RSTB(n7221), .Q(
        \FIFO[64][11] ) );
  DFFARX1 \FIFO_reg[64][10]  ( .D(n2493), .CLK(clk_in), .RSTB(n7221), .Q(
        \FIFO[64][10] ) );
  DFFARX1 \FIFO_reg[64][9]  ( .D(n2492), .CLK(clk_in), .RSTB(n7221), .Q(
        \FIFO[64][9] ) );
  DFFARX1 \FIFO_reg[64][8]  ( .D(n2491), .CLK(clk_in), .RSTB(n7221), .Q(
        \FIFO[64][8] ) );
  DFFARX1 \FIFO_reg[64][7]  ( .D(n2490), .CLK(clk_in), .RSTB(n7221), .Q(
        \FIFO[64][7] ) );
  DFFARX1 \FIFO_reg[64][6]  ( .D(n2489), .CLK(clk_in), .RSTB(n7221), .Q(
        \FIFO[64][6] ) );
  DFFARX1 \FIFO_reg[64][5]  ( .D(n2488), .CLK(clk_in), .RSTB(n7221), .Q(
        \FIFO[64][5] ) );
  DFFARX1 \FIFO_reg[64][4]  ( .D(n2487), .CLK(clk_in), .RSTB(n7221), .Q(
        \FIFO[64][4] ) );
  DFFARX1 \FIFO_reg[64][3]  ( .D(n2486), .CLK(clk_in), .RSTB(n7222), .Q(
        \FIFO[64][3] ) );
  DFFARX1 \FIFO_reg[64][2]  ( .D(n2485), .CLK(clk_in), .RSTB(n7222), .Q(
        \FIFO[64][2] ) );
  DFFARX1 \FIFO_reg[64][1]  ( .D(n2484), .CLK(clk_in), .RSTB(n7222), .Q(
        \FIFO[64][1] ) );
  DFFARX1 \FIFO_reg[64][0]  ( .D(n2483), .CLK(clk_in), .RSTB(n7222), .Q(
        \FIFO[64][0] ) );
  DFFARX1 \FIFO_reg[65][31]  ( .D(n2482), .CLK(clk_in), .RSTB(n7222), .Q(
        \FIFO[65][31] ) );
  DFFARX1 \FIFO_reg[65][30]  ( .D(n2481), .CLK(clk_in), .RSTB(n7222), .Q(
        \FIFO[65][30] ) );
  DFFARX1 \FIFO_reg[65][29]  ( .D(n2480), .CLK(clk_in), .RSTB(n7222), .Q(
        \FIFO[65][29] ) );
  DFFARX1 \FIFO_reg[65][28]  ( .D(n2479), .CLK(clk_in), .RSTB(n7222), .Q(
        \FIFO[65][28] ) );
  DFFARX1 \FIFO_reg[65][27]  ( .D(n2478), .CLK(clk_in), .RSTB(n7222), .Q(
        \FIFO[65][27] ) );
  DFFARX1 \FIFO_reg[65][26]  ( .D(n2477), .CLK(clk_in), .RSTB(n7222), .Q(
        \FIFO[65][26] ) );
  DFFARX1 \FIFO_reg[65][25]  ( .D(n2476), .CLK(clk_in), .RSTB(n7222), .Q(
        \FIFO[65][25] ) );
  DFFARX1 \FIFO_reg[65][24]  ( .D(n2475), .CLK(clk_in), .RSTB(n7222), .Q(
        \FIFO[65][24] ) );
  DFFARX1 \FIFO_reg[65][23]  ( .D(n2474), .CLK(clk_in), .RSTB(n7222), .Q(
        \FIFO[65][23] ) );
  DFFARX1 \FIFO_reg[65][22]  ( .D(n2473), .CLK(clk_in), .RSTB(n7222), .Q(
        \FIFO[65][22] ) );
  DFFARX1 \FIFO_reg[65][21]  ( .D(n2472), .CLK(clk_in), .RSTB(n7222), .Q(
        \FIFO[65][21] ) );
  DFFARX1 \FIFO_reg[65][20]  ( .D(n2471), .CLK(clk_in), .RSTB(n7222), .Q(
        \FIFO[65][20] ) );
  DFFARX1 \FIFO_reg[65][19]  ( .D(n2470), .CLK(clk_in), .RSTB(n7222), .Q(
        \FIFO[65][19] ) );
  DFFARX1 \FIFO_reg[65][18]  ( .D(n2469), .CLK(clk_in), .RSTB(n7222), .Q(
        \FIFO[65][18] ) );
  DFFARX1 \FIFO_reg[65][17]  ( .D(n2468), .CLK(clk_in), .RSTB(n7223), .Q(
        \FIFO[65][17] ) );
  DFFARX1 \FIFO_reg[65][16]  ( .D(n2467), .CLK(clk_in), .RSTB(n7223), .Q(
        \FIFO[65][16] ) );
  DFFARX1 \FIFO_reg[65][15]  ( .D(n2466), .CLK(clk_in), .RSTB(n7223), .Q(
        \FIFO[65][15] ) );
  DFFARX1 \FIFO_reg[65][14]  ( .D(n2465), .CLK(clk_in), .RSTB(n7223), .Q(
        \FIFO[65][14] ) );
  DFFARX1 \FIFO_reg[65][13]  ( .D(n2464), .CLK(clk_in), .RSTB(n7223), .Q(
        \FIFO[65][13] ) );
  DFFARX1 \FIFO_reg[65][12]  ( .D(n2463), .CLK(clk_in), .RSTB(n7223), .Q(
        \FIFO[65][12] ) );
  DFFARX1 \FIFO_reg[65][11]  ( .D(n2462), .CLK(clk_in), .RSTB(n7223), .Q(
        \FIFO[65][11] ) );
  DFFARX1 \FIFO_reg[65][10]  ( .D(n2461), .CLK(clk_in), .RSTB(n7223), .Q(
        \FIFO[65][10] ) );
  DFFARX1 \FIFO_reg[65][9]  ( .D(n2460), .CLK(clk_in), .RSTB(n7223), .Q(
        \FIFO[65][9] ) );
  DFFARX1 \FIFO_reg[65][8]  ( .D(n2459), .CLK(clk_in), .RSTB(n7223), .Q(
        \FIFO[65][8] ) );
  DFFARX1 \FIFO_reg[65][7]  ( .D(n2458), .CLK(clk_in), .RSTB(n7223), .Q(
        \FIFO[65][7] ) );
  DFFARX1 \FIFO_reg[65][6]  ( .D(n2457), .CLK(clk_in), .RSTB(n7223), .Q(
        \FIFO[65][6] ) );
  DFFARX1 \FIFO_reg[65][5]  ( .D(n2456), .CLK(clk_in), .RSTB(n7223), .Q(
        \FIFO[65][5] ) );
  DFFARX1 \FIFO_reg[65][4]  ( .D(n2455), .CLK(clk_in), .RSTB(n7223), .Q(
        \FIFO[65][4] ) );
  DFFARX1 \FIFO_reg[65][3]  ( .D(n2454), .CLK(clk_in), .RSTB(n7223), .Q(
        \FIFO[65][3] ) );
  DFFARX1 \FIFO_reg[65][2]  ( .D(n2453), .CLK(clk_in), .RSTB(n7223), .Q(
        \FIFO[65][2] ) );
  DFFARX1 \FIFO_reg[65][1]  ( .D(n2452), .CLK(clk_in), .RSTB(n7223), .Q(
        \FIFO[65][1] ) );
  DFFARX1 \FIFO_reg[65][0]  ( .D(n2451), .CLK(clk_in), .RSTB(n7223), .Q(
        \FIFO[65][0] ) );
  DFFARX1 \FIFO_reg[66][31]  ( .D(n2450), .CLK(clk_in), .RSTB(n7224), .Q(
        \FIFO[66][31] ) );
  DFFARX1 \FIFO_reg[66][30]  ( .D(n2449), .CLK(clk_in), .RSTB(n7224), .Q(
        \FIFO[66][30] ) );
  DFFARX1 \FIFO_reg[66][29]  ( .D(n2448), .CLK(clk_in), .RSTB(n7224), .Q(
        \FIFO[66][29] ) );
  DFFARX1 \FIFO_reg[66][28]  ( .D(n2447), .CLK(clk_in), .RSTB(n7224), .Q(
        \FIFO[66][28] ) );
  DFFARX1 \FIFO_reg[66][27]  ( .D(n2446), .CLK(clk_in), .RSTB(n7224), .Q(
        \FIFO[66][27] ) );
  DFFARX1 \FIFO_reg[66][26]  ( .D(n2445), .CLK(clk_in), .RSTB(n7224), .Q(
        \FIFO[66][26] ) );
  DFFARX1 \FIFO_reg[66][25]  ( .D(n2444), .CLK(clk_in), .RSTB(n7224), .Q(
        \FIFO[66][25] ) );
  DFFARX1 \FIFO_reg[66][24]  ( .D(n2443), .CLK(clk_in), .RSTB(n7224), .Q(
        \FIFO[66][24] ) );
  DFFARX1 \FIFO_reg[66][23]  ( .D(n2442), .CLK(clk_in), .RSTB(n7224), .Q(
        \FIFO[66][23] ) );
  DFFARX1 \FIFO_reg[66][22]  ( .D(n2441), .CLK(clk_in), .RSTB(n7224), .Q(
        \FIFO[66][22] ) );
  DFFARX1 \FIFO_reg[66][21]  ( .D(n2440), .CLK(clk_in), .RSTB(n7224), .Q(
        \FIFO[66][21] ) );
  DFFARX1 \FIFO_reg[66][20]  ( .D(n2439), .CLK(clk_in), .RSTB(n7224), .Q(
        \FIFO[66][20] ) );
  DFFARX1 \FIFO_reg[66][19]  ( .D(n2438), .CLK(clk_in), .RSTB(n7224), .Q(
        \FIFO[66][19] ) );
  DFFARX1 \FIFO_reg[66][18]  ( .D(n2437), .CLK(clk_in), .RSTB(n7224), .Q(
        \FIFO[66][18] ) );
  DFFARX1 \FIFO_reg[66][17]  ( .D(n2436), .CLK(clk_in), .RSTB(n7224), .Q(
        \FIFO[66][17] ) );
  DFFARX1 \FIFO_reg[66][16]  ( .D(n2435), .CLK(clk_in), .RSTB(n7224), .Q(
        \FIFO[66][16] ) );
  DFFARX1 \FIFO_reg[66][15]  ( .D(n2434), .CLK(clk_in), .RSTB(n7224), .Q(
        \FIFO[66][15] ) );
  DFFARX1 \FIFO_reg[66][14]  ( .D(n2433), .CLK(clk_in), .RSTB(n7224), .Q(
        \FIFO[66][14] ) );
  DFFARX1 \FIFO_reg[66][13]  ( .D(n2432), .CLK(clk_in), .RSTB(n7225), .Q(
        \FIFO[66][13] ) );
  DFFARX1 \FIFO_reg[66][12]  ( .D(n2431), .CLK(clk_in), .RSTB(n7225), .Q(
        \FIFO[66][12] ) );
  DFFARX1 \FIFO_reg[66][11]  ( .D(n2430), .CLK(clk_in), .RSTB(n7225), .Q(
        \FIFO[66][11] ) );
  DFFARX1 \FIFO_reg[66][10]  ( .D(n2429), .CLK(clk_in), .RSTB(n7225), .Q(
        \FIFO[66][10] ) );
  DFFARX1 \FIFO_reg[66][9]  ( .D(n2428), .CLK(clk_in), .RSTB(n7225), .Q(
        \FIFO[66][9] ) );
  DFFARX1 \FIFO_reg[66][8]  ( .D(n2427), .CLK(clk_in), .RSTB(n7225), .Q(
        \FIFO[66][8] ) );
  DFFARX1 \FIFO_reg[66][7]  ( .D(n2426), .CLK(clk_in), .RSTB(n7225), .Q(
        \FIFO[66][7] ) );
  DFFARX1 \FIFO_reg[66][6]  ( .D(n2425), .CLK(clk_in), .RSTB(n7225), .Q(
        \FIFO[66][6] ) );
  DFFARX1 \FIFO_reg[66][5]  ( .D(n2424), .CLK(clk_in), .RSTB(n7225), .Q(
        \FIFO[66][5] ) );
  DFFARX1 \FIFO_reg[66][4]  ( .D(n2423), .CLK(clk_in), .RSTB(n7225), .Q(
        \FIFO[66][4] ) );
  DFFARX1 \FIFO_reg[66][3]  ( .D(n2422), .CLK(clk_in), .RSTB(n7225), .Q(
        \FIFO[66][3] ) );
  DFFARX1 \FIFO_reg[66][2]  ( .D(n2421), .CLK(clk_in), .RSTB(n7225), .Q(
        \FIFO[66][2] ) );
  DFFARX1 \FIFO_reg[66][1]  ( .D(n2420), .CLK(clk_in), .RSTB(n7225), .Q(
        \FIFO[66][1] ) );
  DFFARX1 \FIFO_reg[66][0]  ( .D(n2419), .CLK(clk_in), .RSTB(n7225), .Q(
        \FIFO[66][0] ) );
  DFFARX1 \FIFO_reg[67][31]  ( .D(n2418), .CLK(clk_in), .RSTB(n7225), .Q(
        \FIFO[67][31] ) );
  DFFARX1 \FIFO_reg[67][30]  ( .D(n2417), .CLK(clk_in), .RSTB(n7225), .Q(
        \FIFO[67][30] ) );
  DFFARX1 \FIFO_reg[67][29]  ( .D(n2416), .CLK(clk_in), .RSTB(n7225), .Q(
        \FIFO[67][29] ) );
  DFFARX1 \FIFO_reg[67][28]  ( .D(n2415), .CLK(clk_in), .RSTB(n7225), .Q(
        \FIFO[67][28] ) );
  DFFARX1 \FIFO_reg[67][27]  ( .D(n2414), .CLK(clk_in), .RSTB(n7226), .Q(
        \FIFO[67][27] ) );
  DFFARX1 \FIFO_reg[67][26]  ( .D(n2413), .CLK(clk_in), .RSTB(n7226), .Q(
        \FIFO[67][26] ) );
  DFFARX1 \FIFO_reg[67][25]  ( .D(n2412), .CLK(clk_in), .RSTB(n7226), .Q(
        \FIFO[67][25] ) );
  DFFARX1 \FIFO_reg[67][24]  ( .D(n2411), .CLK(clk_in), .RSTB(n7226), .Q(
        \FIFO[67][24] ) );
  DFFARX1 \FIFO_reg[67][23]  ( .D(n2410), .CLK(clk_in), .RSTB(n7226), .Q(
        \FIFO[67][23] ) );
  DFFARX1 \FIFO_reg[67][22]  ( .D(n2409), .CLK(clk_in), .RSTB(n7226), .Q(
        \FIFO[67][22] ) );
  DFFARX1 \FIFO_reg[67][21]  ( .D(n2408), .CLK(clk_in), .RSTB(n7226), .Q(
        \FIFO[67][21] ) );
  DFFARX1 \FIFO_reg[67][20]  ( .D(n2407), .CLK(clk_in), .RSTB(n7226), .Q(
        \FIFO[67][20] ) );
  DFFARX1 \FIFO_reg[67][19]  ( .D(n2406), .CLK(clk_in), .RSTB(n7226), .Q(
        \FIFO[67][19] ) );
  DFFARX1 \FIFO_reg[67][18]  ( .D(n2405), .CLK(clk_in), .RSTB(n7226), .Q(
        \FIFO[67][18] ) );
  DFFARX1 \FIFO_reg[67][17]  ( .D(n2404), .CLK(clk_in), .RSTB(n7226), .Q(
        \FIFO[67][17] ) );
  DFFARX1 \FIFO_reg[67][16]  ( .D(n2403), .CLK(clk_in), .RSTB(n7226), .Q(
        \FIFO[67][16] ) );
  DFFARX1 \FIFO_reg[67][15]  ( .D(n2402), .CLK(clk_in), .RSTB(n7226), .Q(
        \FIFO[67][15] ) );
  DFFARX1 \FIFO_reg[67][14]  ( .D(n2401), .CLK(clk_in), .RSTB(n7226), .Q(
        \FIFO[67][14] ) );
  DFFARX1 \FIFO_reg[67][13]  ( .D(n2400), .CLK(clk_in), .RSTB(n7226), .Q(
        \FIFO[67][13] ) );
  DFFARX1 \FIFO_reg[67][12]  ( .D(n2399), .CLK(clk_in), .RSTB(n7226), .Q(
        \FIFO[67][12] ) );
  DFFARX1 \FIFO_reg[67][11]  ( .D(n2398), .CLK(clk_in), .RSTB(n7226), .Q(
        \FIFO[67][11] ) );
  DFFARX1 \FIFO_reg[67][10]  ( .D(n2397), .CLK(clk_in), .RSTB(n7226), .Q(
        \FIFO[67][10] ) );
  DFFARX1 \FIFO_reg[67][9]  ( .D(n2396), .CLK(clk_in), .RSTB(n7227), .Q(
        \FIFO[67][9] ) );
  DFFARX1 \FIFO_reg[67][8]  ( .D(n2395), .CLK(clk_in), .RSTB(n7227), .Q(
        \FIFO[67][8] ) );
  DFFARX1 \FIFO_reg[67][7]  ( .D(n2394), .CLK(clk_in), .RSTB(n7227), .Q(
        \FIFO[67][7] ) );
  DFFARX1 \FIFO_reg[67][6]  ( .D(n2393), .CLK(clk_in), .RSTB(n7227), .Q(
        \FIFO[67][6] ) );
  DFFARX1 \FIFO_reg[67][5]  ( .D(n2392), .CLK(clk_in), .RSTB(n7227), .Q(
        \FIFO[67][5] ) );
  DFFARX1 \FIFO_reg[67][4]  ( .D(n2391), .CLK(clk_in), .RSTB(n7227), .Q(
        \FIFO[67][4] ) );
  DFFARX1 \FIFO_reg[67][3]  ( .D(n2390), .CLK(clk_in), .RSTB(n7227), .Q(
        \FIFO[67][3] ) );
  DFFARX1 \FIFO_reg[67][2]  ( .D(n2389), .CLK(clk_in), .RSTB(n7227), .Q(
        \FIFO[67][2] ) );
  DFFARX1 \FIFO_reg[67][1]  ( .D(n2388), .CLK(clk_in), .RSTB(n7227), .Q(
        \FIFO[67][1] ) );
  DFFARX1 \FIFO_reg[67][0]  ( .D(n2387), .CLK(clk_in), .RSTB(n7227), .Q(
        \FIFO[67][0] ) );
  DFFARX1 \FIFO_reg[68][31]  ( .D(n2386), .CLK(clk_in), .RSTB(n7227), .Q(
        \FIFO[68][31] ) );
  DFFARX1 \FIFO_reg[68][30]  ( .D(n2385), .CLK(clk_in), .RSTB(n7227), .Q(
        \FIFO[68][30] ) );
  DFFARX1 \FIFO_reg[68][29]  ( .D(n2384), .CLK(clk_in), .RSTB(n7227), .Q(
        \FIFO[68][29] ) );
  DFFARX1 \FIFO_reg[68][28]  ( .D(n2383), .CLK(clk_in), .RSTB(n7227), .Q(
        \FIFO[68][28] ) );
  DFFARX1 \FIFO_reg[68][27]  ( .D(n2382), .CLK(clk_in), .RSTB(n7227), .Q(
        \FIFO[68][27] ) );
  DFFARX1 \FIFO_reg[68][26]  ( .D(n2381), .CLK(clk_in), .RSTB(n7227), .Q(
        \FIFO[68][26] ) );
  DFFARX1 \FIFO_reg[68][25]  ( .D(n2380), .CLK(clk_in), .RSTB(n7227), .Q(
        \FIFO[68][25] ) );
  DFFARX1 \FIFO_reg[68][24]  ( .D(n2379), .CLK(clk_in), .RSTB(n7227), .Q(
        \FIFO[68][24] ) );
  DFFARX1 \FIFO_reg[68][23]  ( .D(n2378), .CLK(clk_in), .RSTB(n7228), .Q(
        \FIFO[68][23] ) );
  DFFARX1 \FIFO_reg[68][22]  ( .D(n2377), .CLK(clk_in), .RSTB(n7228), .Q(
        \FIFO[68][22] ) );
  DFFARX1 \FIFO_reg[68][21]  ( .D(n2376), .CLK(clk_in), .RSTB(n7228), .Q(
        \FIFO[68][21] ) );
  DFFARX1 \FIFO_reg[68][20]  ( .D(n2375), .CLK(clk_in), .RSTB(n7228), .Q(
        \FIFO[68][20] ) );
  DFFARX1 \FIFO_reg[68][19]  ( .D(n2374), .CLK(clk_in), .RSTB(n7228), .Q(
        \FIFO[68][19] ) );
  DFFARX1 \FIFO_reg[68][18]  ( .D(n2373), .CLK(clk_in), .RSTB(n7228), .Q(
        \FIFO[68][18] ) );
  DFFARX1 \FIFO_reg[68][17]  ( .D(n2372), .CLK(clk_in), .RSTB(n7228), .Q(
        \FIFO[68][17] ) );
  DFFARX1 \FIFO_reg[68][16]  ( .D(n2371), .CLK(clk_in), .RSTB(n7228), .Q(
        \FIFO[68][16] ) );
  DFFARX1 \FIFO_reg[68][15]  ( .D(n2370), .CLK(clk_in), .RSTB(n7228), .Q(
        \FIFO[68][15] ) );
  DFFARX1 \FIFO_reg[68][14]  ( .D(n2369), .CLK(clk_in), .RSTB(n7228), .Q(
        \FIFO[68][14] ) );
  DFFARX1 \FIFO_reg[68][13]  ( .D(n2368), .CLK(clk_in), .RSTB(n7228), .Q(
        \FIFO[68][13] ) );
  DFFARX1 \FIFO_reg[68][12]  ( .D(n2367), .CLK(clk_in), .RSTB(n7228), .Q(
        \FIFO[68][12] ) );
  DFFARX1 \FIFO_reg[68][11]  ( .D(n2366), .CLK(clk_in), .RSTB(n7228), .Q(
        \FIFO[68][11] ) );
  DFFARX1 \FIFO_reg[68][10]  ( .D(n2365), .CLK(clk_in), .RSTB(n7228), .Q(
        \FIFO[68][10] ) );
  DFFARX1 \FIFO_reg[68][9]  ( .D(n2364), .CLK(clk_in), .RSTB(n7228), .Q(
        \FIFO[68][9] ) );
  DFFARX1 \FIFO_reg[68][8]  ( .D(n2363), .CLK(clk_in), .RSTB(n7228), .Q(
        \FIFO[68][8] ) );
  DFFARX1 \FIFO_reg[68][7]  ( .D(n2362), .CLK(clk_in), .RSTB(n7228), .Q(
        \FIFO[68][7] ) );
  DFFARX1 \FIFO_reg[68][6]  ( .D(n2361), .CLK(clk_in), .RSTB(n7228), .Q(
        \FIFO[68][6] ) );
  DFFARX1 \FIFO_reg[68][5]  ( .D(n2360), .CLK(clk_in), .RSTB(n7229), .Q(
        \FIFO[68][5] ) );
  DFFARX1 \FIFO_reg[68][4]  ( .D(n2359), .CLK(clk_in), .RSTB(n7229), .Q(
        \FIFO[68][4] ) );
  DFFARX1 \FIFO_reg[68][3]  ( .D(n2358), .CLK(clk_in), .RSTB(n7229), .Q(
        \FIFO[68][3] ) );
  DFFARX1 \FIFO_reg[68][2]  ( .D(n2357), .CLK(clk_in), .RSTB(n7229), .Q(
        \FIFO[68][2] ) );
  DFFARX1 \FIFO_reg[68][1]  ( .D(n2356), .CLK(clk_in), .RSTB(n7229), .Q(
        \FIFO[68][1] ) );
  DFFARX1 \FIFO_reg[68][0]  ( .D(n2355), .CLK(clk_in), .RSTB(n7229), .Q(
        \FIFO[68][0] ) );
  DFFARX1 \FIFO_reg[69][31]  ( .D(n2354), .CLK(clk_in), .RSTB(n7229), .Q(
        \FIFO[69][31] ) );
  DFFARX1 \FIFO_reg[69][30]  ( .D(n2353), .CLK(clk_in), .RSTB(n7229), .Q(
        \FIFO[69][30] ) );
  DFFARX1 \FIFO_reg[69][29]  ( .D(n2352), .CLK(clk_in), .RSTB(n7229), .Q(
        \FIFO[69][29] ) );
  DFFARX1 \FIFO_reg[69][28]  ( .D(n2351), .CLK(clk_in), .RSTB(n7229), .Q(
        \FIFO[69][28] ) );
  DFFARX1 \FIFO_reg[69][27]  ( .D(n2350), .CLK(clk_in), .RSTB(n7229), .Q(
        \FIFO[69][27] ) );
  DFFARX1 \FIFO_reg[69][26]  ( .D(n2349), .CLK(clk_in), .RSTB(n7229), .Q(
        \FIFO[69][26] ) );
  DFFARX1 \FIFO_reg[69][25]  ( .D(n2348), .CLK(clk_in), .RSTB(n7229), .Q(
        \FIFO[69][25] ) );
  DFFARX1 \FIFO_reg[69][24]  ( .D(n2347), .CLK(clk_in), .RSTB(n7229), .Q(
        \FIFO[69][24] ) );
  DFFARX1 \FIFO_reg[69][23]  ( .D(n2346), .CLK(clk_in), .RSTB(n7229), .Q(
        \FIFO[69][23] ) );
  DFFARX1 \FIFO_reg[69][22]  ( .D(n2345), .CLK(clk_in), .RSTB(n7229), .Q(
        \FIFO[69][22] ) );
  DFFARX1 \FIFO_reg[69][21]  ( .D(n2344), .CLK(clk_in), .RSTB(n7229), .Q(
        \FIFO[69][21] ) );
  DFFARX1 \FIFO_reg[69][20]  ( .D(n2343), .CLK(clk_in), .RSTB(n7229), .Q(
        \FIFO[69][20] ) );
  DFFARX1 \FIFO_reg[69][19]  ( .D(n2342), .CLK(clk_in), .RSTB(n7230), .Q(
        \FIFO[69][19] ) );
  DFFARX1 \FIFO_reg[69][18]  ( .D(n2341), .CLK(clk_in), .RSTB(n7230), .Q(
        \FIFO[69][18] ) );
  DFFARX1 \FIFO_reg[69][17]  ( .D(n2340), .CLK(clk_in), .RSTB(n7230), .Q(
        \FIFO[69][17] ) );
  DFFARX1 \FIFO_reg[69][16]  ( .D(n2339), .CLK(clk_in), .RSTB(n7230), .Q(
        \FIFO[69][16] ) );
  DFFARX1 \FIFO_reg[69][15]  ( .D(n2338), .CLK(clk_in), .RSTB(n7230), .Q(
        \FIFO[69][15] ) );
  DFFARX1 \FIFO_reg[69][14]  ( .D(n2337), .CLK(clk_in), .RSTB(n7230), .Q(
        \FIFO[69][14] ) );
  DFFARX1 \FIFO_reg[69][13]  ( .D(n2336), .CLK(clk_in), .RSTB(n7230), .Q(
        \FIFO[69][13] ) );
  DFFARX1 \FIFO_reg[69][12]  ( .D(n2335), .CLK(clk_in), .RSTB(n7230), .Q(
        \FIFO[69][12] ) );
  DFFARX1 \FIFO_reg[69][11]  ( .D(n2334), .CLK(clk_in), .RSTB(n7230), .Q(
        \FIFO[69][11] ) );
  DFFARX1 \FIFO_reg[69][10]  ( .D(n2333), .CLK(clk_in), .RSTB(n7230), .Q(
        \FIFO[69][10] ) );
  DFFARX1 \FIFO_reg[69][9]  ( .D(n2332), .CLK(clk_in), .RSTB(n7230), .Q(
        \FIFO[69][9] ) );
  DFFARX1 \FIFO_reg[69][8]  ( .D(n2331), .CLK(clk_in), .RSTB(n7230), .Q(
        \FIFO[69][8] ) );
  DFFARX1 \FIFO_reg[69][7]  ( .D(n2330), .CLK(clk_in), .RSTB(n7230), .Q(
        \FIFO[69][7] ) );
  DFFARX1 \FIFO_reg[69][6]  ( .D(n2329), .CLK(clk_in), .RSTB(n7230), .Q(
        \FIFO[69][6] ) );
  DFFARX1 \FIFO_reg[69][5]  ( .D(n2328), .CLK(clk_in), .RSTB(n7230), .Q(
        \FIFO[69][5] ) );
  DFFARX1 \FIFO_reg[69][4]  ( .D(n2327), .CLK(clk_in), .RSTB(n7230), .Q(
        \FIFO[69][4] ) );
  DFFARX1 \FIFO_reg[69][3]  ( .D(n2326), .CLK(clk_in), .RSTB(n7230), .Q(
        \FIFO[69][3] ) );
  DFFARX1 \FIFO_reg[69][2]  ( .D(n2325), .CLK(clk_in), .RSTB(n7230), .Q(
        \FIFO[69][2] ) );
  DFFARX1 \FIFO_reg[69][1]  ( .D(n2324), .CLK(clk_in), .RSTB(n7231), .Q(
        \FIFO[69][1] ) );
  DFFARX1 \FIFO_reg[69][0]  ( .D(n2323), .CLK(clk_in), .RSTB(n7231), .Q(
        \FIFO[69][0] ) );
  DFFARX1 \FIFO_reg[70][31]  ( .D(n2322), .CLK(clk_in), .RSTB(n7231), .Q(
        \FIFO[70][31] ) );
  DFFARX1 \FIFO_reg[70][30]  ( .D(n2321), .CLK(clk_in), .RSTB(n7231), .Q(
        \FIFO[70][30] ) );
  DFFARX1 \FIFO_reg[70][29]  ( .D(n2320), .CLK(clk_in), .RSTB(n7231), .Q(
        \FIFO[70][29] ) );
  DFFARX1 \FIFO_reg[70][28]  ( .D(n2319), .CLK(clk_in), .RSTB(n7231), .Q(
        \FIFO[70][28] ) );
  DFFARX1 \FIFO_reg[70][27]  ( .D(n2318), .CLK(clk_in), .RSTB(n7231), .Q(
        \FIFO[70][27] ) );
  DFFARX1 \FIFO_reg[70][26]  ( .D(n2317), .CLK(clk_in), .RSTB(n7231), .Q(
        \FIFO[70][26] ) );
  DFFARX1 \FIFO_reg[70][25]  ( .D(n2316), .CLK(clk_in), .RSTB(n7231), .Q(
        \FIFO[70][25] ) );
  DFFARX1 \FIFO_reg[70][24]  ( .D(n2315), .CLK(clk_in), .RSTB(n7231), .Q(
        \FIFO[70][24] ) );
  DFFARX1 \FIFO_reg[70][23]  ( .D(n2314), .CLK(clk_in), .RSTB(n7231), .Q(
        \FIFO[70][23] ) );
  DFFARX1 \FIFO_reg[70][22]  ( .D(n2313), .CLK(clk_in), .RSTB(n7231), .Q(
        \FIFO[70][22] ) );
  DFFARX1 \FIFO_reg[70][21]  ( .D(n2312), .CLK(clk_in), .RSTB(n7231), .Q(
        \FIFO[70][21] ) );
  DFFARX1 \FIFO_reg[70][20]  ( .D(n2311), .CLK(clk_in), .RSTB(n7231), .Q(
        \FIFO[70][20] ) );
  DFFARX1 \FIFO_reg[70][19]  ( .D(n2310), .CLK(clk_in), .RSTB(n7231), .Q(
        \FIFO[70][19] ) );
  DFFARX1 \FIFO_reg[70][18]  ( .D(n2309), .CLK(clk_in), .RSTB(n7231), .Q(
        \FIFO[70][18] ) );
  DFFARX1 \FIFO_reg[70][17]  ( .D(n2308), .CLK(clk_in), .RSTB(n7231), .Q(
        \FIFO[70][17] ) );
  DFFARX1 \FIFO_reg[70][16]  ( .D(n2307), .CLK(clk_in), .RSTB(n7231), .Q(
        \FIFO[70][16] ) );
  DFFARX1 \FIFO_reg[70][15]  ( .D(n2306), .CLK(clk_in), .RSTB(n7232), .Q(
        \FIFO[70][15] ) );
  DFFARX1 \FIFO_reg[70][14]  ( .D(n2305), .CLK(clk_in), .RSTB(n7232), .Q(
        \FIFO[70][14] ) );
  DFFARX1 \FIFO_reg[70][13]  ( .D(n2304), .CLK(clk_in), .RSTB(n7232), .Q(
        \FIFO[70][13] ) );
  DFFARX1 \FIFO_reg[70][12]  ( .D(n2303), .CLK(clk_in), .RSTB(n7232), .Q(
        \FIFO[70][12] ) );
  DFFARX1 \FIFO_reg[70][11]  ( .D(n2302), .CLK(clk_in), .RSTB(n7232), .Q(
        \FIFO[70][11] ) );
  DFFARX1 \FIFO_reg[70][10]  ( .D(n2301), .CLK(clk_in), .RSTB(n7232), .Q(
        \FIFO[70][10] ) );
  DFFARX1 \FIFO_reg[70][9]  ( .D(n2300), .CLK(clk_in), .RSTB(n7232), .Q(
        \FIFO[70][9] ) );
  DFFARX1 \FIFO_reg[70][8]  ( .D(n2299), .CLK(clk_in), .RSTB(n7232), .Q(
        \FIFO[70][8] ) );
  DFFARX1 \FIFO_reg[70][7]  ( .D(n2298), .CLK(clk_in), .RSTB(n7232), .Q(
        \FIFO[70][7] ) );
  DFFARX1 \FIFO_reg[70][6]  ( .D(n2297), .CLK(clk_in), .RSTB(n7232), .Q(
        \FIFO[70][6] ) );
  DFFARX1 \FIFO_reg[70][5]  ( .D(n2296), .CLK(clk_in), .RSTB(n7232), .Q(
        \FIFO[70][5] ) );
  DFFARX1 \FIFO_reg[70][4]  ( .D(n2295), .CLK(clk_in), .RSTB(n7232), .Q(
        \FIFO[70][4] ) );
  DFFARX1 \FIFO_reg[70][3]  ( .D(n2294), .CLK(clk_in), .RSTB(n7232), .Q(
        \FIFO[70][3] ) );
  DFFARX1 \FIFO_reg[70][2]  ( .D(n2293), .CLK(clk_in), .RSTB(n7232), .Q(
        \FIFO[70][2] ) );
  DFFARX1 \FIFO_reg[70][1]  ( .D(n2292), .CLK(clk_in), .RSTB(n7232), .Q(
        \FIFO[70][1] ) );
  DFFARX1 \FIFO_reg[70][0]  ( .D(n2291), .CLK(clk_in), .RSTB(n7232), .Q(
        \FIFO[70][0] ) );
  DFFARX1 \FIFO_reg[71][31]  ( .D(n2290), .CLK(clk_in), .RSTB(n7232), .Q(
        \FIFO[71][31] ) );
  DFFARX1 \FIFO_reg[71][30]  ( .D(n2289), .CLK(clk_in), .RSTB(n7232), .Q(
        \FIFO[71][30] ) );
  DFFARX1 \FIFO_reg[71][29]  ( .D(n2288), .CLK(clk_in), .RSTB(n7233), .Q(
        \FIFO[71][29] ) );
  DFFARX1 \FIFO_reg[71][28]  ( .D(n2287), .CLK(clk_in), .RSTB(n7233), .Q(
        \FIFO[71][28] ) );
  DFFARX1 \FIFO_reg[71][27]  ( .D(n2286), .CLK(clk_in), .RSTB(n7233), .Q(
        \FIFO[71][27] ) );
  DFFARX1 \FIFO_reg[71][26]  ( .D(n2285), .CLK(clk_in), .RSTB(n7233), .Q(
        \FIFO[71][26] ) );
  DFFARX1 \FIFO_reg[71][25]  ( .D(n2284), .CLK(clk_in), .RSTB(n7233), .Q(
        \FIFO[71][25] ) );
  DFFARX1 \FIFO_reg[71][24]  ( .D(n2283), .CLK(clk_in), .RSTB(n7233), .Q(
        \FIFO[71][24] ) );
  DFFARX1 \FIFO_reg[71][23]  ( .D(n2282), .CLK(clk_in), .RSTB(n7233), .Q(
        \FIFO[71][23] ) );
  DFFARX1 \FIFO_reg[71][22]  ( .D(n2281), .CLK(clk_in), .RSTB(n7233), .Q(
        \FIFO[71][22] ) );
  DFFARX1 \FIFO_reg[71][21]  ( .D(n2280), .CLK(clk_in), .RSTB(n7233), .Q(
        \FIFO[71][21] ) );
  DFFARX1 \FIFO_reg[71][20]  ( .D(n2279), .CLK(clk_in), .RSTB(n7233), .Q(
        \FIFO[71][20] ) );
  DFFARX1 \FIFO_reg[71][19]  ( .D(n2278), .CLK(clk_in), .RSTB(n7233), .Q(
        \FIFO[71][19] ) );
  DFFARX1 \FIFO_reg[71][18]  ( .D(n2277), .CLK(clk_in), .RSTB(n7233), .Q(
        \FIFO[71][18] ) );
  DFFARX1 \FIFO_reg[71][17]  ( .D(n2276), .CLK(clk_in), .RSTB(n7233), .Q(
        \FIFO[71][17] ) );
  DFFARX1 \FIFO_reg[71][16]  ( .D(n2275), .CLK(clk_in), .RSTB(n7233), .Q(
        \FIFO[71][16] ) );
  DFFARX1 \FIFO_reg[71][15]  ( .D(n2274), .CLK(clk_in), .RSTB(n7233), .Q(
        \FIFO[71][15] ) );
  DFFARX1 \FIFO_reg[71][14]  ( .D(n2273), .CLK(clk_in), .RSTB(n7233), .Q(
        \FIFO[71][14] ) );
  DFFARX1 \FIFO_reg[71][13]  ( .D(n2272), .CLK(clk_in), .RSTB(n7233), .Q(
        \FIFO[71][13] ) );
  DFFARX1 \FIFO_reg[71][12]  ( .D(n2271), .CLK(clk_in), .RSTB(n7233), .Q(
        \FIFO[71][12] ) );
  DFFARX1 \FIFO_reg[71][11]  ( .D(n2270), .CLK(clk_in), .RSTB(n7234), .Q(
        \FIFO[71][11] ) );
  DFFARX1 \FIFO_reg[71][10]  ( .D(n2269), .CLK(clk_in), .RSTB(n7234), .Q(
        \FIFO[71][10] ) );
  DFFARX1 \FIFO_reg[71][9]  ( .D(n2268), .CLK(clk_in), .RSTB(n7234), .Q(
        \FIFO[71][9] ) );
  DFFARX1 \FIFO_reg[71][8]  ( .D(n2267), .CLK(clk_in), .RSTB(n7234), .Q(
        \FIFO[71][8] ) );
  DFFARX1 \FIFO_reg[71][7]  ( .D(n2266), .CLK(clk_in), .RSTB(n7234), .Q(
        \FIFO[71][7] ) );
  DFFARX1 \FIFO_reg[71][6]  ( .D(n2265), .CLK(clk_in), .RSTB(n7234), .Q(
        \FIFO[71][6] ) );
  DFFARX1 \FIFO_reg[71][5]  ( .D(n2264), .CLK(clk_in), .RSTB(n7234), .Q(
        \FIFO[71][5] ) );
  DFFARX1 \FIFO_reg[71][4]  ( .D(n2263), .CLK(clk_in), .RSTB(n7234), .Q(
        \FIFO[71][4] ) );
  DFFARX1 \FIFO_reg[71][3]  ( .D(n2262), .CLK(clk_in), .RSTB(n7234), .Q(
        \FIFO[71][3] ) );
  DFFARX1 \FIFO_reg[71][2]  ( .D(n2261), .CLK(clk_in), .RSTB(n7234), .Q(
        \FIFO[71][2] ) );
  DFFARX1 \FIFO_reg[71][1]  ( .D(n2260), .CLK(clk_in), .RSTB(n7234), .Q(
        \FIFO[71][1] ) );
  DFFARX1 \FIFO_reg[71][0]  ( .D(n2259), .CLK(clk_in), .RSTB(n7234), .Q(
        \FIFO[71][0] ) );
  DFFARX1 \FIFO_reg[72][31]  ( .D(n2258), .CLK(clk_in), .RSTB(n7234), .Q(
        \FIFO[72][31] ) );
  DFFARX1 \FIFO_reg[72][30]  ( .D(n2257), .CLK(clk_in), .RSTB(n7234), .Q(
        \FIFO[72][30] ) );
  DFFARX1 \FIFO_reg[72][29]  ( .D(n2256), .CLK(clk_in), .RSTB(n7234), .Q(
        \FIFO[72][29] ) );
  DFFARX1 \FIFO_reg[72][28]  ( .D(n2255), .CLK(clk_in), .RSTB(n7234), .Q(
        \FIFO[72][28] ) );
  DFFARX1 \FIFO_reg[72][27]  ( .D(n2254), .CLK(clk_in), .RSTB(n7234), .Q(
        \FIFO[72][27] ) );
  DFFARX1 \FIFO_reg[72][26]  ( .D(n2253), .CLK(clk_in), .RSTB(n7234), .Q(
        \FIFO[72][26] ) );
  DFFARX1 \FIFO_reg[72][25]  ( .D(n2252), .CLK(clk_in), .RSTB(n7235), .Q(
        \FIFO[72][25] ) );
  DFFARX1 \FIFO_reg[72][24]  ( .D(n2251), .CLK(clk_in), .RSTB(n7235), .Q(
        \FIFO[72][24] ) );
  DFFARX1 \FIFO_reg[72][23]  ( .D(n2250), .CLK(clk_in), .RSTB(n7235), .Q(
        \FIFO[72][23] ) );
  DFFARX1 \FIFO_reg[72][22]  ( .D(n2249), .CLK(clk_in), .RSTB(n7235), .Q(
        \FIFO[72][22] ) );
  DFFARX1 \FIFO_reg[72][21]  ( .D(n2248), .CLK(clk_in), .RSTB(n7235), .Q(
        \FIFO[72][21] ) );
  DFFARX1 \FIFO_reg[72][20]  ( .D(n2247), .CLK(clk_in), .RSTB(n7235), .Q(
        \FIFO[72][20] ) );
  DFFARX1 \FIFO_reg[72][19]  ( .D(n2246), .CLK(clk_in), .RSTB(n7235), .Q(
        \FIFO[72][19] ) );
  DFFARX1 \FIFO_reg[72][18]  ( .D(n2245), .CLK(clk_in), .RSTB(n7235), .Q(
        \FIFO[72][18] ) );
  DFFARX1 \FIFO_reg[72][17]  ( .D(n2244), .CLK(clk_in), .RSTB(n7235), .Q(
        \FIFO[72][17] ) );
  DFFARX1 \FIFO_reg[72][16]  ( .D(n2243), .CLK(clk_in), .RSTB(n7235), .Q(
        \FIFO[72][16] ) );
  DFFARX1 \FIFO_reg[72][15]  ( .D(n2242), .CLK(clk_in), .RSTB(n7235), .Q(
        \FIFO[72][15] ) );
  DFFARX1 \FIFO_reg[72][14]  ( .D(n2241), .CLK(clk_in), .RSTB(n7235), .Q(
        \FIFO[72][14] ) );
  DFFARX1 \FIFO_reg[72][13]  ( .D(n2240), .CLK(clk_in), .RSTB(n7235), .Q(
        \FIFO[72][13] ) );
  DFFARX1 \FIFO_reg[72][12]  ( .D(n2239), .CLK(clk_in), .RSTB(n7235), .Q(
        \FIFO[72][12] ) );
  DFFARX1 \FIFO_reg[72][11]  ( .D(n2238), .CLK(clk_in), .RSTB(n7235), .Q(
        \FIFO[72][11] ) );
  DFFARX1 \FIFO_reg[72][10]  ( .D(n2237), .CLK(clk_in), .RSTB(n7235), .Q(
        \FIFO[72][10] ) );
  DFFARX1 \FIFO_reg[72][9]  ( .D(n2236), .CLK(clk_in), .RSTB(n7235), .Q(
        \FIFO[72][9] ) );
  DFFARX1 \FIFO_reg[72][8]  ( .D(n2235), .CLK(clk_in), .RSTB(n7235), .Q(
        \FIFO[72][8] ) );
  DFFARX1 \FIFO_reg[72][7]  ( .D(n2234), .CLK(clk_in), .RSTB(n7236), .Q(
        \FIFO[72][7] ) );
  DFFARX1 \FIFO_reg[72][6]  ( .D(n2233), .CLK(clk_in), .RSTB(n7236), .Q(
        \FIFO[72][6] ) );
  DFFARX1 \FIFO_reg[72][5]  ( .D(n2232), .CLK(clk_in), .RSTB(n7236), .Q(
        \FIFO[72][5] ) );
  DFFARX1 \FIFO_reg[72][4]  ( .D(n2231), .CLK(clk_in), .RSTB(n7236), .Q(
        \FIFO[72][4] ) );
  DFFARX1 \FIFO_reg[72][3]  ( .D(n2230), .CLK(clk_in), .RSTB(n7236), .Q(
        \FIFO[72][3] ) );
  DFFARX1 \FIFO_reg[72][2]  ( .D(n2229), .CLK(clk_in), .RSTB(n7236), .Q(
        \FIFO[72][2] ) );
  DFFARX1 \FIFO_reg[72][1]  ( .D(n2228), .CLK(clk_in), .RSTB(n7236), .Q(
        \FIFO[72][1] ) );
  DFFARX1 \FIFO_reg[72][0]  ( .D(n2227), .CLK(clk_in), .RSTB(n7236), .Q(
        \FIFO[72][0] ) );
  DFFARX1 \FIFO_reg[73][31]  ( .D(n2226), .CLK(clk_in), .RSTB(n7236), .Q(
        \FIFO[73][31] ) );
  DFFARX1 \FIFO_reg[73][30]  ( .D(n2225), .CLK(clk_in), .RSTB(n7236), .Q(
        \FIFO[73][30] ) );
  DFFARX1 \FIFO_reg[73][29]  ( .D(n2224), .CLK(clk_in), .RSTB(n7236), .Q(
        \FIFO[73][29] ) );
  DFFARX1 \FIFO_reg[73][28]  ( .D(n2223), .CLK(clk_in), .RSTB(n7236), .Q(
        \FIFO[73][28] ) );
  DFFARX1 \FIFO_reg[73][27]  ( .D(n2222), .CLK(clk_in), .RSTB(n7236), .Q(
        \FIFO[73][27] ) );
  DFFARX1 \FIFO_reg[73][26]  ( .D(n2221), .CLK(clk_in), .RSTB(n7236), .Q(
        \FIFO[73][26] ) );
  DFFARX1 \FIFO_reg[73][25]  ( .D(n2220), .CLK(clk_in), .RSTB(n7236), .Q(
        \FIFO[73][25] ) );
  DFFARX1 \FIFO_reg[73][24]  ( .D(n2219), .CLK(clk_in), .RSTB(n7236), .Q(
        \FIFO[73][24] ) );
  DFFARX1 \FIFO_reg[73][23]  ( .D(n2218), .CLK(clk_in), .RSTB(n7236), .Q(
        \FIFO[73][23] ) );
  DFFARX1 \FIFO_reg[73][22]  ( .D(n2217), .CLK(clk_in), .RSTB(n7236), .Q(
        \FIFO[73][22] ) );
  DFFARX1 \FIFO_reg[73][21]  ( .D(n2216), .CLK(clk_in), .RSTB(n7237), .Q(
        \FIFO[73][21] ) );
  DFFARX1 \FIFO_reg[73][20]  ( .D(n2215), .CLK(clk_in), .RSTB(n7237), .Q(
        \FIFO[73][20] ) );
  DFFARX1 \FIFO_reg[73][19]  ( .D(n2214), .CLK(clk_in), .RSTB(n7237), .Q(
        \FIFO[73][19] ) );
  DFFARX1 \FIFO_reg[73][18]  ( .D(n2213), .CLK(clk_in), .RSTB(n7237), .Q(
        \FIFO[73][18] ) );
  DFFARX1 \FIFO_reg[73][17]  ( .D(n2212), .CLK(clk_in), .RSTB(n7237), .Q(
        \FIFO[73][17] ) );
  DFFARX1 \FIFO_reg[73][16]  ( .D(n2211), .CLK(clk_in), .RSTB(n7237), .Q(
        \FIFO[73][16] ) );
  DFFARX1 \FIFO_reg[73][15]  ( .D(n2210), .CLK(clk_in), .RSTB(n7237), .Q(
        \FIFO[73][15] ) );
  DFFARX1 \FIFO_reg[73][14]  ( .D(n2209), .CLK(clk_in), .RSTB(n7237), .Q(
        \FIFO[73][14] ) );
  DFFARX1 \FIFO_reg[73][13]  ( .D(n2208), .CLK(clk_in), .RSTB(n7237), .Q(
        \FIFO[73][13] ) );
  DFFARX1 \FIFO_reg[73][12]  ( .D(n2207), .CLK(clk_in), .RSTB(n7237), .Q(
        \FIFO[73][12] ) );
  DFFARX1 \FIFO_reg[73][11]  ( .D(n2206), .CLK(clk_in), .RSTB(n7237), .Q(
        \FIFO[73][11] ) );
  DFFARX1 \FIFO_reg[73][10]  ( .D(n2205), .CLK(clk_in), .RSTB(n7237), .Q(
        \FIFO[73][10] ) );
  DFFARX1 \FIFO_reg[73][9]  ( .D(n2204), .CLK(clk_in), .RSTB(n7237), .Q(
        \FIFO[73][9] ) );
  DFFARX1 \FIFO_reg[73][8]  ( .D(n2203), .CLK(clk_in), .RSTB(n7237), .Q(
        \FIFO[73][8] ) );
  DFFARX1 \FIFO_reg[73][7]  ( .D(n2202), .CLK(clk_in), .RSTB(n7237), .Q(
        \FIFO[73][7] ) );
  DFFARX1 \FIFO_reg[73][6]  ( .D(n2201), .CLK(clk_in), .RSTB(n7237), .Q(
        \FIFO[73][6] ) );
  DFFARX1 \FIFO_reg[73][5]  ( .D(n2200), .CLK(clk_in), .RSTB(n7237), .Q(
        \FIFO[73][5] ) );
  DFFARX1 \FIFO_reg[73][4]  ( .D(n2199), .CLK(clk_in), .RSTB(n7237), .Q(
        \FIFO[73][4] ) );
  DFFARX1 \FIFO_reg[73][3]  ( .D(n2198), .CLK(clk_in), .RSTB(n7238), .Q(
        \FIFO[73][3] ) );
  DFFARX1 \FIFO_reg[73][2]  ( .D(n2197), .CLK(clk_in), .RSTB(n7238), .Q(
        \FIFO[73][2] ) );
  DFFARX1 \FIFO_reg[73][1]  ( .D(n2196), .CLK(clk_in), .RSTB(n7238), .Q(
        \FIFO[73][1] ) );
  DFFARX1 \FIFO_reg[73][0]  ( .D(n2195), .CLK(clk_in), .RSTB(n7238), .Q(
        \FIFO[73][0] ) );
  DFFARX1 \FIFO_reg[74][31]  ( .D(n2194), .CLK(clk_in), .RSTB(n7238), .Q(
        \FIFO[74][31] ) );
  DFFARX1 \FIFO_reg[74][30]  ( .D(n2193), .CLK(clk_in), .RSTB(n7238), .Q(
        \FIFO[74][30] ) );
  DFFARX1 \FIFO_reg[74][29]  ( .D(n2192), .CLK(clk_in), .RSTB(n7238), .Q(
        \FIFO[74][29] ) );
  DFFARX1 \FIFO_reg[74][28]  ( .D(n2191), .CLK(clk_in), .RSTB(n7238), .Q(
        \FIFO[74][28] ) );
  DFFARX1 \FIFO_reg[74][27]  ( .D(n2190), .CLK(clk_in), .RSTB(n7238), .Q(
        \FIFO[74][27] ) );
  DFFARX1 \FIFO_reg[74][26]  ( .D(n2189), .CLK(clk_in), .RSTB(n7238), .Q(
        \FIFO[74][26] ) );
  DFFARX1 \FIFO_reg[74][25]  ( .D(n2188), .CLK(clk_in), .RSTB(n7238), .Q(
        \FIFO[74][25] ) );
  DFFARX1 \FIFO_reg[74][24]  ( .D(n2187), .CLK(clk_in), .RSTB(n7238), .Q(
        \FIFO[74][24] ) );
  DFFARX1 \FIFO_reg[74][23]  ( .D(n2186), .CLK(clk_in), .RSTB(n7238), .Q(
        \FIFO[74][23] ) );
  DFFARX1 \FIFO_reg[74][22]  ( .D(n2185), .CLK(clk_in), .RSTB(n7238), .Q(
        \FIFO[74][22] ) );
  DFFARX1 \FIFO_reg[74][21]  ( .D(n2184), .CLK(clk_in), .RSTB(n7238), .Q(
        \FIFO[74][21] ) );
  DFFARX1 \FIFO_reg[74][20]  ( .D(n2183), .CLK(clk_in), .RSTB(n7238), .Q(
        \FIFO[74][20] ) );
  DFFARX1 \FIFO_reg[74][19]  ( .D(n2182), .CLK(clk_in), .RSTB(n7238), .Q(
        \FIFO[74][19] ) );
  DFFARX1 \FIFO_reg[74][18]  ( .D(n2181), .CLK(clk_in), .RSTB(n7238), .Q(
        \FIFO[74][18] ) );
  DFFARX1 \FIFO_reg[74][17]  ( .D(n2180), .CLK(clk_in), .RSTB(n7239), .Q(
        \FIFO[74][17] ) );
  DFFARX1 \FIFO_reg[74][16]  ( .D(n2179), .CLK(clk_in), .RSTB(n7239), .Q(
        \FIFO[74][16] ) );
  DFFARX1 \FIFO_reg[74][15]  ( .D(n2178), .CLK(clk_in), .RSTB(n7239), .Q(
        \FIFO[74][15] ) );
  DFFARX1 \FIFO_reg[74][14]  ( .D(n2177), .CLK(clk_in), .RSTB(n7239), .Q(
        \FIFO[74][14] ) );
  DFFARX1 \FIFO_reg[74][13]  ( .D(n2176), .CLK(clk_in), .RSTB(n7239), .Q(
        \FIFO[74][13] ) );
  DFFARX1 \FIFO_reg[74][12]  ( .D(n2175), .CLK(clk_in), .RSTB(n7239), .Q(
        \FIFO[74][12] ) );
  DFFARX1 \FIFO_reg[74][11]  ( .D(n2174), .CLK(clk_in), .RSTB(n7239), .Q(
        \FIFO[74][11] ) );
  DFFARX1 \FIFO_reg[74][10]  ( .D(n2173), .CLK(clk_in), .RSTB(n7239), .Q(
        \FIFO[74][10] ) );
  DFFARX1 \FIFO_reg[74][9]  ( .D(n2172), .CLK(clk_in), .RSTB(n7239), .Q(
        \FIFO[74][9] ) );
  DFFARX1 \FIFO_reg[74][8]  ( .D(n2171), .CLK(clk_in), .RSTB(n7239), .Q(
        \FIFO[74][8] ) );
  DFFARX1 \FIFO_reg[74][7]  ( .D(n2170), .CLK(clk_in), .RSTB(n7239), .Q(
        \FIFO[74][7] ) );
  DFFARX1 \FIFO_reg[74][6]  ( .D(n2169), .CLK(clk_in), .RSTB(n7239), .Q(
        \FIFO[74][6] ) );
  DFFARX1 \FIFO_reg[74][5]  ( .D(n2168), .CLK(clk_in), .RSTB(n7239), .Q(
        \FIFO[74][5] ) );
  DFFARX1 \FIFO_reg[74][4]  ( .D(n2167), .CLK(clk_in), .RSTB(n7239), .Q(
        \FIFO[74][4] ) );
  DFFARX1 \FIFO_reg[74][3]  ( .D(n2166), .CLK(clk_in), .RSTB(n7239), .Q(
        \FIFO[74][3] ) );
  DFFARX1 \FIFO_reg[74][2]  ( .D(n2165), .CLK(clk_in), .RSTB(n7239), .Q(
        \FIFO[74][2] ) );
  DFFARX1 \FIFO_reg[74][1]  ( .D(n2164), .CLK(clk_in), .RSTB(n7239), .Q(
        \FIFO[74][1] ) );
  DFFARX1 \FIFO_reg[74][0]  ( .D(n2163), .CLK(clk_in), .RSTB(n7239), .Q(
        \FIFO[74][0] ) );
  DFFARX1 \FIFO_reg[75][31]  ( .D(n2162), .CLK(clk_in), .RSTB(n7240), .Q(
        \FIFO[75][31] ) );
  DFFARX1 \FIFO_reg[75][30]  ( .D(n2161), .CLK(clk_in), .RSTB(n7240), .Q(
        \FIFO[75][30] ) );
  DFFARX1 \FIFO_reg[75][29]  ( .D(n2160), .CLK(clk_in), .RSTB(n7240), .Q(
        \FIFO[75][29] ) );
  DFFARX1 \FIFO_reg[75][28]  ( .D(n2159), .CLK(clk_in), .RSTB(n7240), .Q(
        \FIFO[75][28] ) );
  DFFARX1 \FIFO_reg[75][27]  ( .D(n2158), .CLK(clk_in), .RSTB(n7240), .Q(
        \FIFO[75][27] ) );
  DFFARX1 \FIFO_reg[75][26]  ( .D(n2157), .CLK(clk_in), .RSTB(n7240), .Q(
        \FIFO[75][26] ) );
  DFFARX1 \FIFO_reg[75][25]  ( .D(n2156), .CLK(clk_in), .RSTB(n7240), .Q(
        \FIFO[75][25] ) );
  DFFARX1 \FIFO_reg[75][24]  ( .D(n2155), .CLK(clk_in), .RSTB(n7240), .Q(
        \FIFO[75][24] ) );
  DFFARX1 \FIFO_reg[75][23]  ( .D(n2154), .CLK(clk_in), .RSTB(n7240), .Q(
        \FIFO[75][23] ) );
  DFFARX1 \FIFO_reg[75][22]  ( .D(n2153), .CLK(clk_in), .RSTB(n7240), .Q(
        \FIFO[75][22] ) );
  DFFARX1 \FIFO_reg[75][21]  ( .D(n2152), .CLK(clk_in), .RSTB(n7240), .Q(
        \FIFO[75][21] ) );
  DFFARX1 \FIFO_reg[75][20]  ( .D(n2151), .CLK(clk_in), .RSTB(n7240), .Q(
        \FIFO[75][20] ) );
  DFFARX1 \FIFO_reg[75][19]  ( .D(n2150), .CLK(clk_in), .RSTB(n7240), .Q(
        \FIFO[75][19] ) );
  DFFARX1 \FIFO_reg[75][18]  ( .D(n2149), .CLK(clk_in), .RSTB(n7240), .Q(
        \FIFO[75][18] ) );
  DFFARX1 \FIFO_reg[75][17]  ( .D(n2148), .CLK(clk_in), .RSTB(n7240), .Q(
        \FIFO[75][17] ) );
  DFFARX1 \FIFO_reg[75][16]  ( .D(n2147), .CLK(clk_in), .RSTB(n7240), .Q(
        \FIFO[75][16] ) );
  DFFARX1 \FIFO_reg[75][15]  ( .D(n2146), .CLK(clk_in), .RSTB(n7240), .Q(
        \FIFO[75][15] ) );
  DFFARX1 \FIFO_reg[75][14]  ( .D(n2145), .CLK(clk_in), .RSTB(n7240), .Q(
        \FIFO[75][14] ) );
  DFFARX1 \FIFO_reg[75][13]  ( .D(n2144), .CLK(clk_in), .RSTB(n7241), .Q(
        \FIFO[75][13] ) );
  DFFARX1 \FIFO_reg[75][12]  ( .D(n2143), .CLK(clk_in), .RSTB(n7241), .Q(
        \FIFO[75][12] ) );
  DFFARX1 \FIFO_reg[75][11]  ( .D(n2142), .CLK(clk_in), .RSTB(n7241), .Q(
        \FIFO[75][11] ) );
  DFFARX1 \FIFO_reg[75][10]  ( .D(n2141), .CLK(clk_in), .RSTB(n7241), .Q(
        \FIFO[75][10] ) );
  DFFARX1 \FIFO_reg[75][9]  ( .D(n2140), .CLK(clk_in), .RSTB(n7241), .Q(
        \FIFO[75][9] ) );
  DFFARX1 \FIFO_reg[75][8]  ( .D(n2139), .CLK(clk_in), .RSTB(n7241), .Q(
        \FIFO[75][8] ) );
  DFFARX1 \FIFO_reg[75][7]  ( .D(n2138), .CLK(clk_in), .RSTB(n7241), .Q(
        \FIFO[75][7] ) );
  DFFARX1 \FIFO_reg[75][6]  ( .D(n2137), .CLK(clk_in), .RSTB(n7241), .Q(
        \FIFO[75][6] ) );
  DFFARX1 \FIFO_reg[75][5]  ( .D(n2136), .CLK(clk_in), .RSTB(n7241), .Q(
        \FIFO[75][5] ) );
  DFFARX1 \FIFO_reg[75][4]  ( .D(n2135), .CLK(clk_in), .RSTB(n7241), .Q(
        \FIFO[75][4] ) );
  DFFARX1 \FIFO_reg[75][3]  ( .D(n2134), .CLK(clk_in), .RSTB(n7241), .Q(
        \FIFO[75][3] ) );
  DFFARX1 \FIFO_reg[75][2]  ( .D(n2133), .CLK(clk_in), .RSTB(n7241), .Q(
        \FIFO[75][2] ) );
  DFFARX1 \FIFO_reg[75][1]  ( .D(n2132), .CLK(clk_in), .RSTB(n7241), .Q(
        \FIFO[75][1] ) );
  DFFARX1 \FIFO_reg[75][0]  ( .D(n2131), .CLK(clk_in), .RSTB(n7241), .Q(
        \FIFO[75][0] ) );
  DFFARX1 \FIFO_reg[76][31]  ( .D(n2130), .CLK(clk_in), .RSTB(n7241), .Q(
        \FIFO[76][31] ) );
  DFFARX1 \FIFO_reg[76][30]  ( .D(n2129), .CLK(clk_in), .RSTB(n7241), .Q(
        \FIFO[76][30] ) );
  DFFARX1 \FIFO_reg[76][29]  ( .D(n2128), .CLK(clk_in), .RSTB(n7241), .Q(
        \FIFO[76][29] ) );
  DFFARX1 \FIFO_reg[76][28]  ( .D(n2127), .CLK(clk_in), .RSTB(n7241), .Q(
        \FIFO[76][28] ) );
  DFFARX1 \FIFO_reg[76][27]  ( .D(n2126), .CLK(clk_in), .RSTB(n7242), .Q(
        \FIFO[76][27] ) );
  DFFARX1 \FIFO_reg[76][26]  ( .D(n2125), .CLK(clk_in), .RSTB(n7242), .Q(
        \FIFO[76][26] ) );
  DFFARX1 \FIFO_reg[76][25]  ( .D(n2124), .CLK(clk_in), .RSTB(n7242), .Q(
        \FIFO[76][25] ) );
  DFFARX1 \FIFO_reg[76][24]  ( .D(n2123), .CLK(clk_in), .RSTB(n7242), .Q(
        \FIFO[76][24] ) );
  DFFARX1 \FIFO_reg[76][23]  ( .D(n2122), .CLK(clk_in), .RSTB(n7242), .Q(
        \FIFO[76][23] ) );
  DFFARX1 \FIFO_reg[76][22]  ( .D(n2121), .CLK(clk_in), .RSTB(n7242), .Q(
        \FIFO[76][22] ) );
  DFFARX1 \FIFO_reg[76][21]  ( .D(n2120), .CLK(clk_in), .RSTB(n7242), .Q(
        \FIFO[76][21] ) );
  DFFARX1 \FIFO_reg[76][20]  ( .D(n2119), .CLK(clk_in), .RSTB(n7242), .Q(
        \FIFO[76][20] ) );
  DFFARX1 \FIFO_reg[76][19]  ( .D(n2118), .CLK(clk_in), .RSTB(n7242), .Q(
        \FIFO[76][19] ) );
  DFFARX1 \FIFO_reg[76][18]  ( .D(n2117), .CLK(clk_in), .RSTB(n7242), .Q(
        \FIFO[76][18] ) );
  DFFARX1 \FIFO_reg[76][17]  ( .D(n2116), .CLK(clk_in), .RSTB(n7242), .Q(
        \FIFO[76][17] ) );
  DFFARX1 \FIFO_reg[76][16]  ( .D(n2115), .CLK(clk_in), .RSTB(n7242), .Q(
        \FIFO[76][16] ) );
  DFFARX1 \FIFO_reg[76][15]  ( .D(n2114), .CLK(clk_in), .RSTB(n7242), .Q(
        \FIFO[76][15] ) );
  DFFARX1 \FIFO_reg[76][14]  ( .D(n2113), .CLK(clk_in), .RSTB(n7242), .Q(
        \FIFO[76][14] ) );
  DFFARX1 \FIFO_reg[76][13]  ( .D(n2112), .CLK(clk_in), .RSTB(n7242), .Q(
        \FIFO[76][13] ) );
  DFFARX1 \FIFO_reg[76][12]  ( .D(n2111), .CLK(clk_in), .RSTB(n7242), .Q(
        \FIFO[76][12] ) );
  DFFARX1 \FIFO_reg[76][11]  ( .D(n2110), .CLK(clk_in), .RSTB(n7242), .Q(
        \FIFO[76][11] ) );
  DFFARX1 \FIFO_reg[76][10]  ( .D(n2109), .CLK(clk_in), .RSTB(n7242), .Q(
        \FIFO[76][10] ) );
  DFFARX1 \FIFO_reg[76][9]  ( .D(n2108), .CLK(clk_in), .RSTB(n7243), .Q(
        \FIFO[76][9] ) );
  DFFARX1 \FIFO_reg[76][8]  ( .D(n2107), .CLK(clk_in), .RSTB(n7243), .Q(
        \FIFO[76][8] ) );
  DFFARX1 \FIFO_reg[76][7]  ( .D(n2106), .CLK(clk_in), .RSTB(n7243), .Q(
        \FIFO[76][7] ) );
  DFFARX1 \FIFO_reg[76][6]  ( .D(n2105), .CLK(clk_in), .RSTB(n7243), .Q(
        \FIFO[76][6] ) );
  DFFARX1 \FIFO_reg[76][5]  ( .D(n2104), .CLK(clk_in), .RSTB(n7243), .Q(
        \FIFO[76][5] ) );
  DFFARX1 \FIFO_reg[76][4]  ( .D(n2103), .CLK(clk_in), .RSTB(n7243), .Q(
        \FIFO[76][4] ) );
  DFFARX1 \FIFO_reg[76][3]  ( .D(n2102), .CLK(clk_in), .RSTB(n7243), .Q(
        \FIFO[76][3] ) );
  DFFARX1 \FIFO_reg[76][2]  ( .D(n2101), .CLK(clk_in), .RSTB(n7243), .Q(
        \FIFO[76][2] ) );
  DFFARX1 \FIFO_reg[76][1]  ( .D(n2100), .CLK(clk_in), .RSTB(n7243), .Q(
        \FIFO[76][1] ) );
  DFFARX1 \FIFO_reg[76][0]  ( .D(n2099), .CLK(clk_in), .RSTB(n7243), .Q(
        \FIFO[76][0] ) );
  DFFARX1 \FIFO_reg[77][31]  ( .D(n2098), .CLK(clk_in), .RSTB(n7243), .Q(
        \FIFO[77][31] ) );
  DFFARX1 \FIFO_reg[77][30]  ( .D(n2097), .CLK(clk_in), .RSTB(n7243), .Q(
        \FIFO[77][30] ) );
  DFFARX1 \FIFO_reg[77][29]  ( .D(n2096), .CLK(clk_in), .RSTB(n7243), .Q(
        \FIFO[77][29] ) );
  DFFARX1 \FIFO_reg[77][28]  ( .D(n2095), .CLK(clk_in), .RSTB(n7243), .Q(
        \FIFO[77][28] ) );
  DFFARX1 \FIFO_reg[77][27]  ( .D(n2094), .CLK(clk_in), .RSTB(n7243), .Q(
        \FIFO[77][27] ) );
  DFFARX1 \FIFO_reg[77][26]  ( .D(n2093), .CLK(clk_in), .RSTB(n7243), .Q(
        \FIFO[77][26] ) );
  DFFARX1 \FIFO_reg[77][25]  ( .D(n2092), .CLK(clk_in), .RSTB(n7243), .Q(
        \FIFO[77][25] ) );
  DFFARX1 \FIFO_reg[77][24]  ( .D(n2091), .CLK(clk_in), .RSTB(n7243), .Q(
        \FIFO[77][24] ) );
  DFFARX1 \FIFO_reg[77][23]  ( .D(n2090), .CLK(clk_in), .RSTB(n7244), .Q(
        \FIFO[77][23] ) );
  DFFARX1 \FIFO_reg[77][22]  ( .D(n2089), .CLK(clk_in), .RSTB(n7244), .Q(
        \FIFO[77][22] ) );
  DFFARX1 \FIFO_reg[77][21]  ( .D(n2088), .CLK(clk_in), .RSTB(n7244), .Q(
        \FIFO[77][21] ) );
  DFFARX1 \FIFO_reg[77][20]  ( .D(n2087), .CLK(clk_in), .RSTB(n7244), .Q(
        \FIFO[77][20] ) );
  DFFARX1 \FIFO_reg[77][19]  ( .D(n2086), .CLK(clk_in), .RSTB(n7244), .Q(
        \FIFO[77][19] ) );
  DFFARX1 \FIFO_reg[77][18]  ( .D(n2085), .CLK(clk_in), .RSTB(n7244), .Q(
        \FIFO[77][18] ) );
  DFFARX1 \FIFO_reg[77][17]  ( .D(n2084), .CLK(clk_in), .RSTB(n7244), .Q(
        \FIFO[77][17] ) );
  DFFARX1 \FIFO_reg[77][16]  ( .D(n2083), .CLK(clk_in), .RSTB(n7244), .Q(
        \FIFO[77][16] ) );
  DFFARX1 \FIFO_reg[77][15]  ( .D(n2082), .CLK(clk_in), .RSTB(n7244), .Q(
        \FIFO[77][15] ) );
  DFFARX1 \FIFO_reg[77][14]  ( .D(n2081), .CLK(clk_in), .RSTB(n7244), .Q(
        \FIFO[77][14] ) );
  DFFARX1 \FIFO_reg[77][13]  ( .D(n2080), .CLK(clk_in), .RSTB(n7244), .Q(
        \FIFO[77][13] ) );
  DFFARX1 \FIFO_reg[77][12]  ( .D(n2079), .CLK(clk_in), .RSTB(n7244), .Q(
        \FIFO[77][12] ) );
  DFFARX1 \FIFO_reg[77][11]  ( .D(n2078), .CLK(clk_in), .RSTB(n7244), .Q(
        \FIFO[77][11] ) );
  DFFARX1 \FIFO_reg[77][10]  ( .D(n2077), .CLK(clk_in), .RSTB(n7244), .Q(
        \FIFO[77][10] ) );
  DFFARX1 \FIFO_reg[77][9]  ( .D(n2076), .CLK(clk_in), .RSTB(n7244), .Q(
        \FIFO[77][9] ) );
  DFFARX1 \FIFO_reg[77][8]  ( .D(n2075), .CLK(clk_in), .RSTB(n7244), .Q(
        \FIFO[77][8] ) );
  DFFARX1 \FIFO_reg[77][7]  ( .D(n2074), .CLK(clk_in), .RSTB(n7244), .Q(
        \FIFO[77][7] ) );
  DFFARX1 \FIFO_reg[77][6]  ( .D(n2073), .CLK(clk_in), .RSTB(n7244), .Q(
        \FIFO[77][6] ) );
  DFFARX1 \FIFO_reg[77][5]  ( .D(n2072), .CLK(clk_in), .RSTB(n7245), .Q(
        \FIFO[77][5] ) );
  DFFARX1 \FIFO_reg[77][4]  ( .D(n2071), .CLK(clk_in), .RSTB(n7245), .Q(
        \FIFO[77][4] ) );
  DFFARX1 \FIFO_reg[77][3]  ( .D(n2070), .CLK(clk_in), .RSTB(n7245), .Q(
        \FIFO[77][3] ) );
  DFFARX1 \FIFO_reg[77][2]  ( .D(n2069), .CLK(clk_in), .RSTB(n7245), .Q(
        \FIFO[77][2] ) );
  DFFARX1 \FIFO_reg[77][1]  ( .D(n2068), .CLK(clk_in), .RSTB(n7245), .Q(
        \FIFO[77][1] ) );
  DFFARX1 \FIFO_reg[77][0]  ( .D(n2067), .CLK(clk_in), .RSTB(n7245), .Q(
        \FIFO[77][0] ) );
  DFFARX1 \FIFO_reg[78][31]  ( .D(n2066), .CLK(clk_in), .RSTB(n7245), .Q(
        \FIFO[78][31] ) );
  DFFARX1 \FIFO_reg[78][30]  ( .D(n2065), .CLK(clk_in), .RSTB(n7245), .Q(
        \FIFO[78][30] ) );
  DFFARX1 \FIFO_reg[78][29]  ( .D(n2064), .CLK(clk_in), .RSTB(n7245), .Q(
        \FIFO[78][29] ) );
  DFFARX1 \FIFO_reg[78][28]  ( .D(n2063), .CLK(clk_in), .RSTB(n7245), .Q(
        \FIFO[78][28] ) );
  DFFARX1 \FIFO_reg[78][27]  ( .D(n2062), .CLK(clk_in), .RSTB(n7245), .Q(
        \FIFO[78][27] ) );
  DFFARX1 \FIFO_reg[78][26]  ( .D(n2061), .CLK(clk_in), .RSTB(n7245), .Q(
        \FIFO[78][26] ) );
  DFFARX1 \FIFO_reg[78][25]  ( .D(n2060), .CLK(clk_in), .RSTB(n7245), .Q(
        \FIFO[78][25] ) );
  DFFARX1 \FIFO_reg[78][24]  ( .D(n2059), .CLK(clk_in), .RSTB(n7245), .Q(
        \FIFO[78][24] ) );
  DFFARX1 \FIFO_reg[78][23]  ( .D(n2058), .CLK(clk_in), .RSTB(n7245), .Q(
        \FIFO[78][23] ) );
  DFFARX1 \FIFO_reg[78][22]  ( .D(n2057), .CLK(clk_in), .RSTB(n7245), .Q(
        \FIFO[78][22] ) );
  DFFARX1 \FIFO_reg[78][21]  ( .D(n2056), .CLK(clk_in), .RSTB(n7245), .Q(
        \FIFO[78][21] ) );
  DFFARX1 \FIFO_reg[78][20]  ( .D(n2055), .CLK(clk_in), .RSTB(n7245), .Q(
        \FIFO[78][20] ) );
  DFFARX1 \FIFO_reg[78][19]  ( .D(n2054), .CLK(clk_in), .RSTB(n7246), .Q(
        \FIFO[78][19] ) );
  DFFARX1 \FIFO_reg[78][18]  ( .D(n2053), .CLK(clk_in), .RSTB(n7246), .Q(
        \FIFO[78][18] ) );
  DFFARX1 \FIFO_reg[78][17]  ( .D(n2052), .CLK(clk_in), .RSTB(n7246), .Q(
        \FIFO[78][17] ) );
  DFFARX1 \FIFO_reg[78][16]  ( .D(n2051), .CLK(clk_in), .RSTB(n7246), .Q(
        \FIFO[78][16] ) );
  DFFARX1 \FIFO_reg[78][15]  ( .D(n2050), .CLK(clk_in), .RSTB(n7246), .Q(
        \FIFO[78][15] ) );
  DFFARX1 \FIFO_reg[78][14]  ( .D(n2049), .CLK(clk_in), .RSTB(n7246), .Q(
        \FIFO[78][14] ) );
  DFFARX1 \FIFO_reg[78][13]  ( .D(n2048), .CLK(clk_in), .RSTB(n7246), .Q(
        \FIFO[78][13] ) );
  DFFARX1 \FIFO_reg[78][12]  ( .D(n2047), .CLK(clk_in), .RSTB(n7246), .Q(
        \FIFO[78][12] ) );
  DFFARX1 \FIFO_reg[78][11]  ( .D(n2046), .CLK(clk_in), .RSTB(n7246), .Q(
        \FIFO[78][11] ) );
  DFFARX1 \FIFO_reg[78][10]  ( .D(n2045), .CLK(clk_in), .RSTB(n7246), .Q(
        \FIFO[78][10] ) );
  DFFARX1 \FIFO_reg[78][9]  ( .D(n2044), .CLK(clk_in), .RSTB(n7246), .Q(
        \FIFO[78][9] ) );
  DFFARX1 \FIFO_reg[78][8]  ( .D(n2043), .CLK(clk_in), .RSTB(n7246), .Q(
        \FIFO[78][8] ) );
  DFFARX1 \FIFO_reg[78][7]  ( .D(n2042), .CLK(clk_in), .RSTB(n7246), .Q(
        \FIFO[78][7] ) );
  DFFARX1 \FIFO_reg[78][6]  ( .D(n2041), .CLK(clk_in), .RSTB(n7246), .Q(
        \FIFO[78][6] ) );
  DFFARX1 \FIFO_reg[78][5]  ( .D(n2040), .CLK(clk_in), .RSTB(n7246), .Q(
        \FIFO[78][5] ) );
  DFFARX1 \FIFO_reg[78][4]  ( .D(n2039), .CLK(clk_in), .RSTB(n7246), .Q(
        \FIFO[78][4] ) );
  DFFARX1 \FIFO_reg[78][3]  ( .D(n2038), .CLK(clk_in), .RSTB(n7246), .Q(
        \FIFO[78][3] ) );
  DFFARX1 \FIFO_reg[78][2]  ( .D(n2037), .CLK(clk_in), .RSTB(n7246), .Q(
        \FIFO[78][2] ) );
  DFFARX1 \FIFO_reg[78][1]  ( .D(n2036), .CLK(clk_in), .RSTB(n7247), .Q(
        \FIFO[78][1] ) );
  DFFARX1 \FIFO_reg[78][0]  ( .D(n2035), .CLK(clk_in), .RSTB(n7247), .Q(
        \FIFO[78][0] ) );
  DFFARX1 \FIFO_reg[79][31]  ( .D(n2034), .CLK(clk_in), .RSTB(n7247), .Q(
        \FIFO[79][31] ) );
  DFFARX1 \FIFO_reg[79][30]  ( .D(n2033), .CLK(clk_in), .RSTB(n7247), .Q(
        \FIFO[79][30] ) );
  DFFARX1 \FIFO_reg[79][29]  ( .D(n2032), .CLK(clk_in), .RSTB(n7247), .Q(
        \FIFO[79][29] ) );
  DFFARX1 \FIFO_reg[79][28]  ( .D(n2031), .CLK(clk_in), .RSTB(n7247), .Q(
        \FIFO[79][28] ) );
  DFFARX1 \FIFO_reg[79][27]  ( .D(n2030), .CLK(clk_in), .RSTB(n7247), .Q(
        \FIFO[79][27] ) );
  DFFARX1 \FIFO_reg[79][26]  ( .D(n2029), .CLK(clk_in), .RSTB(n7247), .Q(
        \FIFO[79][26] ) );
  DFFARX1 \FIFO_reg[79][25]  ( .D(n2028), .CLK(clk_in), .RSTB(n7247), .Q(
        \FIFO[79][25] ) );
  DFFARX1 \FIFO_reg[79][24]  ( .D(n2027), .CLK(clk_in), .RSTB(n7247), .Q(
        \FIFO[79][24] ) );
  DFFARX1 \FIFO_reg[79][23]  ( .D(n2026), .CLK(clk_in), .RSTB(n7247), .Q(
        \FIFO[79][23] ) );
  DFFARX1 \FIFO_reg[79][22]  ( .D(n2025), .CLK(clk_in), .RSTB(n7247), .Q(
        \FIFO[79][22] ) );
  DFFARX1 \FIFO_reg[79][21]  ( .D(n2024), .CLK(clk_in), .RSTB(n7247), .Q(
        \FIFO[79][21] ) );
  DFFARX1 \FIFO_reg[79][20]  ( .D(n2023), .CLK(clk_in), .RSTB(n7247), .Q(
        \FIFO[79][20] ) );
  DFFARX1 \FIFO_reg[79][19]  ( .D(n2022), .CLK(clk_in), .RSTB(n7247), .Q(
        \FIFO[79][19] ) );
  DFFARX1 \FIFO_reg[79][18]  ( .D(n2021), .CLK(clk_in), .RSTB(n7247), .Q(
        \FIFO[79][18] ) );
  DFFARX1 \FIFO_reg[79][17]  ( .D(n2020), .CLK(clk_in), .RSTB(n7247), .Q(
        \FIFO[79][17] ) );
  DFFARX1 \FIFO_reg[79][16]  ( .D(n2019), .CLK(clk_in), .RSTB(n7247), .Q(
        \FIFO[79][16] ) );
  DFFARX1 \FIFO_reg[79][15]  ( .D(n2018), .CLK(clk_in), .RSTB(n7248), .Q(
        \FIFO[79][15] ) );
  DFFARX1 \FIFO_reg[79][14]  ( .D(n2017), .CLK(clk_in), .RSTB(n7248), .Q(
        \FIFO[79][14] ) );
  DFFARX1 \FIFO_reg[79][13]  ( .D(n2016), .CLK(clk_in), .RSTB(n7248), .Q(
        \FIFO[79][13] ) );
  DFFARX1 \FIFO_reg[79][12]  ( .D(n2015), .CLK(clk_in), .RSTB(n7248), .Q(
        \FIFO[79][12] ) );
  DFFARX1 \FIFO_reg[79][11]  ( .D(n2014), .CLK(clk_in), .RSTB(n7248), .Q(
        \FIFO[79][11] ) );
  DFFARX1 \FIFO_reg[79][10]  ( .D(n2013), .CLK(clk_in), .RSTB(n7248), .Q(
        \FIFO[79][10] ) );
  DFFARX1 \FIFO_reg[79][9]  ( .D(n2012), .CLK(clk_in), .RSTB(n7248), .Q(
        \FIFO[79][9] ) );
  DFFARX1 \FIFO_reg[79][8]  ( .D(n2011), .CLK(clk_in), .RSTB(n7248), .Q(
        \FIFO[79][8] ) );
  DFFARX1 \FIFO_reg[79][7]  ( .D(n2010), .CLK(clk_in), .RSTB(n7248), .Q(
        \FIFO[79][7] ) );
  DFFARX1 \FIFO_reg[79][6]  ( .D(n2009), .CLK(clk_in), .RSTB(n7248), .Q(
        \FIFO[79][6] ) );
  DFFARX1 \FIFO_reg[79][5]  ( .D(n2008), .CLK(clk_in), .RSTB(n7248), .Q(
        \FIFO[79][5] ) );
  DFFARX1 \FIFO_reg[79][4]  ( .D(n2007), .CLK(clk_in), .RSTB(n7248), .Q(
        \FIFO[79][4] ) );
  DFFARX1 \FIFO_reg[79][3]  ( .D(n2006), .CLK(clk_in), .RSTB(n7248), .Q(
        \FIFO[79][3] ) );
  DFFARX1 \FIFO_reg[79][2]  ( .D(n2005), .CLK(clk_in), .RSTB(n7248), .Q(
        \FIFO[79][2] ) );
  DFFARX1 \FIFO_reg[79][1]  ( .D(n2004), .CLK(clk_in), .RSTB(n7248), .Q(
        \FIFO[79][1] ) );
  DFFARX1 \FIFO_reg[79][0]  ( .D(n2003), .CLK(clk_in), .RSTB(n7248), .Q(
        \FIFO[79][0] ) );
  DFFARX1 \FIFO_reg[80][31]  ( .D(n2002), .CLK(clk_in), .RSTB(n7248), .Q(
        \FIFO[80][31] ) );
  DFFARX1 \FIFO_reg[80][30]  ( .D(n2001), .CLK(clk_in), .RSTB(n7248), .Q(
        \FIFO[80][30] ) );
  DFFARX1 \FIFO_reg[80][29]  ( .D(n2000), .CLK(clk_in), .RSTB(n7249), .Q(
        \FIFO[80][29] ) );
  DFFARX1 \FIFO_reg[80][28]  ( .D(n1999), .CLK(clk_in), .RSTB(n7249), .Q(
        \FIFO[80][28] ) );
  DFFARX1 \FIFO_reg[80][27]  ( .D(n1998), .CLK(clk_in), .RSTB(n7249), .Q(
        \FIFO[80][27] ) );
  DFFARX1 \FIFO_reg[80][26]  ( .D(n1997), .CLK(clk_in), .RSTB(n7249), .Q(
        \FIFO[80][26] ) );
  DFFARX1 \FIFO_reg[80][25]  ( .D(n1996), .CLK(clk_in), .RSTB(n7249), .Q(
        \FIFO[80][25] ) );
  DFFARX1 \FIFO_reg[80][24]  ( .D(n1995), .CLK(clk_in), .RSTB(n7249), .Q(
        \FIFO[80][24] ) );
  DFFARX1 \FIFO_reg[80][23]  ( .D(n1994), .CLK(clk_in), .RSTB(n7249), .Q(
        \FIFO[80][23] ) );
  DFFARX1 \FIFO_reg[80][22]  ( .D(n1993), .CLK(clk_in), .RSTB(n7249), .Q(
        \FIFO[80][22] ) );
  DFFARX1 \FIFO_reg[80][21]  ( .D(n1992), .CLK(clk_in), .RSTB(n7249), .Q(
        \FIFO[80][21] ) );
  DFFARX1 \FIFO_reg[80][20]  ( .D(n1991), .CLK(clk_in), .RSTB(n7249), .Q(
        \FIFO[80][20] ) );
  DFFARX1 \FIFO_reg[80][19]  ( .D(n1990), .CLK(clk_in), .RSTB(n7249), .Q(
        \FIFO[80][19] ) );
  DFFARX1 \FIFO_reg[80][18]  ( .D(n1989), .CLK(clk_in), .RSTB(n7249), .Q(
        \FIFO[80][18] ) );
  DFFARX1 \FIFO_reg[80][17]  ( .D(n1988), .CLK(clk_in), .RSTB(n7249), .Q(
        \FIFO[80][17] ) );
  DFFARX1 \FIFO_reg[80][16]  ( .D(n1987), .CLK(clk_in), .RSTB(n7249), .Q(
        \FIFO[80][16] ) );
  DFFARX1 \FIFO_reg[80][15]  ( .D(n1986), .CLK(clk_in), .RSTB(n7249), .Q(
        \FIFO[80][15] ) );
  DFFARX1 \FIFO_reg[80][14]  ( .D(n1985), .CLK(clk_in), .RSTB(n7249), .Q(
        \FIFO[80][14] ) );
  DFFARX1 \FIFO_reg[80][13]  ( .D(n1984), .CLK(clk_in), .RSTB(n7249), .Q(
        \FIFO[80][13] ) );
  DFFARX1 \FIFO_reg[80][12]  ( .D(n1983), .CLK(clk_in), .RSTB(n7249), .Q(
        \FIFO[80][12] ) );
  DFFARX1 \FIFO_reg[80][11]  ( .D(n1982), .CLK(clk_in), .RSTB(n7250), .Q(
        \FIFO[80][11] ) );
  DFFARX1 \FIFO_reg[80][10]  ( .D(n1981), .CLK(clk_in), .RSTB(n7250), .Q(
        \FIFO[80][10] ) );
  DFFARX1 \FIFO_reg[80][9]  ( .D(n1980), .CLK(clk_in), .RSTB(n7250), .Q(
        \FIFO[80][9] ) );
  DFFARX1 \FIFO_reg[80][8]  ( .D(n1979), .CLK(clk_in), .RSTB(n7250), .Q(
        \FIFO[80][8] ) );
  DFFARX1 \FIFO_reg[80][7]  ( .D(n1978), .CLK(clk_in), .RSTB(n7250), .Q(
        \FIFO[80][7] ) );
  DFFARX1 \FIFO_reg[80][6]  ( .D(n1977), .CLK(clk_in), .RSTB(n7250), .Q(
        \FIFO[80][6] ) );
  DFFARX1 \FIFO_reg[80][5]  ( .D(n1976), .CLK(clk_in), .RSTB(n7250), .Q(
        \FIFO[80][5] ) );
  DFFARX1 \FIFO_reg[80][4]  ( .D(n1975), .CLK(clk_in), .RSTB(n7250), .Q(
        \FIFO[80][4] ) );
  DFFARX1 \FIFO_reg[80][3]  ( .D(n1974), .CLK(clk_in), .RSTB(n7250), .Q(
        \FIFO[80][3] ) );
  DFFARX1 \FIFO_reg[80][2]  ( .D(n1973), .CLK(clk_in), .RSTB(n7250), .Q(
        \FIFO[80][2] ) );
  DFFARX1 \FIFO_reg[80][1]  ( .D(n1972), .CLK(clk_in), .RSTB(n7250), .Q(
        \FIFO[80][1] ) );
  DFFARX1 \FIFO_reg[80][0]  ( .D(n1971), .CLK(clk_in), .RSTB(n7250), .Q(
        \FIFO[80][0] ) );
  DFFARX1 \FIFO_reg[81][31]  ( .D(n1970), .CLK(clk_in), .RSTB(n7250), .Q(
        \FIFO[81][31] ) );
  DFFARX1 \FIFO_reg[81][30]  ( .D(n1969), .CLK(clk_in), .RSTB(n7250), .Q(
        \FIFO[81][30] ) );
  DFFARX1 \FIFO_reg[81][29]  ( .D(n1968), .CLK(clk_in), .RSTB(n7250), .Q(
        \FIFO[81][29] ) );
  DFFARX1 \FIFO_reg[81][28]  ( .D(n1967), .CLK(clk_in), .RSTB(n7250), .Q(
        \FIFO[81][28] ) );
  DFFARX1 \FIFO_reg[81][27]  ( .D(n1966), .CLK(clk_in), .RSTB(n7250), .Q(
        \FIFO[81][27] ) );
  DFFARX1 \FIFO_reg[81][26]  ( .D(n1965), .CLK(clk_in), .RSTB(n7250), .Q(
        \FIFO[81][26] ) );
  DFFARX1 \FIFO_reg[81][25]  ( .D(n1964), .CLK(clk_in), .RSTB(n7251), .Q(
        \FIFO[81][25] ) );
  DFFARX1 \FIFO_reg[81][24]  ( .D(n1963), .CLK(clk_in), .RSTB(n7251), .Q(
        \FIFO[81][24] ) );
  DFFARX1 \FIFO_reg[81][23]  ( .D(n1962), .CLK(clk_in), .RSTB(n7251), .Q(
        \FIFO[81][23] ) );
  DFFARX1 \FIFO_reg[81][22]  ( .D(n1961), .CLK(clk_in), .RSTB(n7251), .Q(
        \FIFO[81][22] ) );
  DFFARX1 \FIFO_reg[81][21]  ( .D(n1960), .CLK(clk_in), .RSTB(n7251), .Q(
        \FIFO[81][21] ) );
  DFFARX1 \FIFO_reg[81][20]  ( .D(n1959), .CLK(clk_in), .RSTB(n7251), .Q(
        \FIFO[81][20] ) );
  DFFARX1 \FIFO_reg[81][19]  ( .D(n1958), .CLK(clk_in), .RSTB(n7251), .Q(
        \FIFO[81][19] ) );
  DFFARX1 \FIFO_reg[81][18]  ( .D(n1957), .CLK(clk_in), .RSTB(n7251), .Q(
        \FIFO[81][18] ) );
  DFFARX1 \FIFO_reg[81][17]  ( .D(n1956), .CLK(clk_in), .RSTB(n7251), .Q(
        \FIFO[81][17] ) );
  DFFARX1 \FIFO_reg[81][16]  ( .D(n1955), .CLK(clk_in), .RSTB(n7251), .Q(
        \FIFO[81][16] ) );
  DFFARX1 \FIFO_reg[81][15]  ( .D(n1954), .CLK(clk_in), .RSTB(n7251), .Q(
        \FIFO[81][15] ) );
  DFFARX1 \FIFO_reg[81][14]  ( .D(n1953), .CLK(clk_in), .RSTB(n7251), .Q(
        \FIFO[81][14] ) );
  DFFARX1 \FIFO_reg[81][13]  ( .D(n1952), .CLK(clk_in), .RSTB(n7251), .Q(
        \FIFO[81][13] ) );
  DFFARX1 \FIFO_reg[81][12]  ( .D(n1951), .CLK(clk_in), .RSTB(n7251), .Q(
        \FIFO[81][12] ) );
  DFFARX1 \FIFO_reg[81][11]  ( .D(n1950), .CLK(clk_in), .RSTB(n7251), .Q(
        \FIFO[81][11] ) );
  DFFARX1 \FIFO_reg[81][10]  ( .D(n1949), .CLK(clk_in), .RSTB(n7251), .Q(
        \FIFO[81][10] ) );
  DFFARX1 \FIFO_reg[81][9]  ( .D(n1948), .CLK(clk_in), .RSTB(n7251), .Q(
        \FIFO[81][9] ) );
  DFFARX1 \FIFO_reg[81][8]  ( .D(n1947), .CLK(clk_in), .RSTB(n7251), .Q(
        \FIFO[81][8] ) );
  DFFARX1 \FIFO_reg[81][7]  ( .D(n1946), .CLK(clk_in), .RSTB(n7252), .Q(
        \FIFO[81][7] ) );
  DFFARX1 \FIFO_reg[81][6]  ( .D(n1945), .CLK(clk_in), .RSTB(n7252), .Q(
        \FIFO[81][6] ) );
  DFFARX1 \FIFO_reg[81][5]  ( .D(n1944), .CLK(clk_in), .RSTB(n7252), .Q(
        \FIFO[81][5] ) );
  DFFARX1 \FIFO_reg[81][4]  ( .D(n1943), .CLK(clk_in), .RSTB(n7252), .Q(
        \FIFO[81][4] ) );
  DFFARX1 \FIFO_reg[81][3]  ( .D(n1942), .CLK(clk_in), .RSTB(n7252), .Q(
        \FIFO[81][3] ) );
  DFFARX1 \FIFO_reg[81][2]  ( .D(n1941), .CLK(clk_in), .RSTB(n7252), .Q(
        \FIFO[81][2] ) );
  DFFARX1 \FIFO_reg[81][1]  ( .D(n1940), .CLK(clk_in), .RSTB(n7252), .Q(
        \FIFO[81][1] ) );
  DFFARX1 \FIFO_reg[81][0]  ( .D(n1939), .CLK(clk_in), .RSTB(n7252), .Q(
        \FIFO[81][0] ) );
  DFFARX1 \FIFO_reg[82][31]  ( .D(n1938), .CLK(clk_in), .RSTB(n7252), .Q(
        \FIFO[82][31] ) );
  DFFARX1 \FIFO_reg[82][30]  ( .D(n1937), .CLK(clk_in), .RSTB(n7252), .Q(
        \FIFO[82][30] ) );
  DFFARX1 \FIFO_reg[82][29]  ( .D(n1936), .CLK(clk_in), .RSTB(n7252), .Q(
        \FIFO[82][29] ) );
  DFFARX1 \FIFO_reg[82][28]  ( .D(n1935), .CLK(clk_in), .RSTB(n7252), .Q(
        \FIFO[82][28] ) );
  DFFARX1 \FIFO_reg[82][27]  ( .D(n1934), .CLK(clk_in), .RSTB(n7252), .Q(
        \FIFO[82][27] ) );
  DFFARX1 \FIFO_reg[82][26]  ( .D(n1933), .CLK(clk_in), .RSTB(n7252), .Q(
        \FIFO[82][26] ) );
  DFFARX1 \FIFO_reg[82][25]  ( .D(n1932), .CLK(clk_in), .RSTB(n7252), .Q(
        \FIFO[82][25] ) );
  DFFARX1 \FIFO_reg[82][24]  ( .D(n1931), .CLK(clk_in), .RSTB(n7252), .Q(
        \FIFO[82][24] ) );
  DFFARX1 \FIFO_reg[82][23]  ( .D(n1930), .CLK(clk_in), .RSTB(n7252), .Q(
        \FIFO[82][23] ) );
  DFFARX1 \FIFO_reg[82][22]  ( .D(n1929), .CLK(clk_in), .RSTB(n7252), .Q(
        \FIFO[82][22] ) );
  DFFARX1 \FIFO_reg[82][21]  ( .D(n1928), .CLK(clk_in), .RSTB(n7253), .Q(
        \FIFO[82][21] ) );
  DFFARX1 \FIFO_reg[82][20]  ( .D(n1927), .CLK(clk_in), .RSTB(n7253), .Q(
        \FIFO[82][20] ) );
  DFFARX1 \FIFO_reg[82][19]  ( .D(n1926), .CLK(clk_in), .RSTB(n7253), .Q(
        \FIFO[82][19] ) );
  DFFARX1 \FIFO_reg[82][18]  ( .D(n1925), .CLK(clk_in), .RSTB(n7253), .Q(
        \FIFO[82][18] ) );
  DFFARX1 \FIFO_reg[82][17]  ( .D(n1924), .CLK(clk_in), .RSTB(n7253), .Q(
        \FIFO[82][17] ) );
  DFFARX1 \FIFO_reg[82][16]  ( .D(n1923), .CLK(clk_in), .RSTB(n7253), .Q(
        \FIFO[82][16] ) );
  DFFARX1 \FIFO_reg[82][15]  ( .D(n1922), .CLK(clk_in), .RSTB(n7253), .Q(
        \FIFO[82][15] ) );
  DFFARX1 \FIFO_reg[82][14]  ( .D(n1921), .CLK(clk_in), .RSTB(n7253), .Q(
        \FIFO[82][14] ) );
  DFFARX1 \FIFO_reg[82][13]  ( .D(n1920), .CLK(clk_in), .RSTB(n7253), .Q(
        \FIFO[82][13] ) );
  DFFARX1 \FIFO_reg[82][12]  ( .D(n1919), .CLK(clk_in), .RSTB(n7253), .Q(
        \FIFO[82][12] ) );
  DFFARX1 \FIFO_reg[82][11]  ( .D(n1918), .CLK(clk_in), .RSTB(n7253), .Q(
        \FIFO[82][11] ) );
  DFFARX1 \FIFO_reg[82][10]  ( .D(n1917), .CLK(clk_in), .RSTB(n7253), .Q(
        \FIFO[82][10] ) );
  DFFARX1 \FIFO_reg[82][9]  ( .D(n1916), .CLK(clk_in), .RSTB(n7253), .Q(
        \FIFO[82][9] ) );
  DFFARX1 \FIFO_reg[82][8]  ( .D(n1915), .CLK(clk_in), .RSTB(n7253), .Q(
        \FIFO[82][8] ) );
  DFFARX1 \FIFO_reg[82][7]  ( .D(n1914), .CLK(clk_in), .RSTB(n7253), .Q(
        \FIFO[82][7] ) );
  DFFARX1 \FIFO_reg[82][6]  ( .D(n1913), .CLK(clk_in), .RSTB(n7253), .Q(
        \FIFO[82][6] ) );
  DFFARX1 \FIFO_reg[82][5]  ( .D(n1912), .CLK(clk_in), .RSTB(n7253), .Q(
        \FIFO[82][5] ) );
  DFFARX1 \FIFO_reg[82][4]  ( .D(n1911), .CLK(clk_in), .RSTB(n7253), .Q(
        \FIFO[82][4] ) );
  DFFARX1 \FIFO_reg[82][3]  ( .D(n1910), .CLK(clk_in), .RSTB(n7254), .Q(
        \FIFO[82][3] ) );
  DFFARX1 \FIFO_reg[82][2]  ( .D(n1909), .CLK(clk_in), .RSTB(n7254), .Q(
        \FIFO[82][2] ) );
  DFFARX1 \FIFO_reg[82][1]  ( .D(n1908), .CLK(clk_in), .RSTB(n7254), .Q(
        \FIFO[82][1] ) );
  DFFARX1 \FIFO_reg[82][0]  ( .D(n1907), .CLK(clk_in), .RSTB(n7254), .Q(
        \FIFO[82][0] ) );
  DFFARX1 \FIFO_reg[83][31]  ( .D(n1906), .CLK(clk_in), .RSTB(n7254), .Q(
        \FIFO[83][31] ) );
  DFFARX1 \FIFO_reg[83][30]  ( .D(n1905), .CLK(clk_in), .RSTB(n7254), .Q(
        \FIFO[83][30] ) );
  DFFARX1 \FIFO_reg[83][29]  ( .D(n1904), .CLK(clk_in), .RSTB(n7254), .Q(
        \FIFO[83][29] ) );
  DFFARX1 \FIFO_reg[83][28]  ( .D(n1903), .CLK(clk_in), .RSTB(n7254), .Q(
        \FIFO[83][28] ) );
  DFFARX1 \FIFO_reg[83][27]  ( .D(n1902), .CLK(clk_in), .RSTB(n7254), .Q(
        \FIFO[83][27] ) );
  DFFARX1 \FIFO_reg[83][26]  ( .D(n1901), .CLK(clk_in), .RSTB(n7254), .Q(
        \FIFO[83][26] ) );
  DFFARX1 \FIFO_reg[83][25]  ( .D(n1900), .CLK(clk_in), .RSTB(n7254), .Q(
        \FIFO[83][25] ) );
  DFFARX1 \FIFO_reg[83][24]  ( .D(n1899), .CLK(clk_in), .RSTB(n7254), .Q(
        \FIFO[83][24] ) );
  DFFARX1 \FIFO_reg[83][23]  ( .D(n1898), .CLK(clk_in), .RSTB(n7254), .Q(
        \FIFO[83][23] ) );
  DFFARX1 \FIFO_reg[83][22]  ( .D(n1897), .CLK(clk_in), .RSTB(n7254), .Q(
        \FIFO[83][22] ) );
  DFFARX1 \FIFO_reg[83][21]  ( .D(n1896), .CLK(clk_in), .RSTB(n7254), .Q(
        \FIFO[83][21] ) );
  DFFARX1 \FIFO_reg[83][20]  ( .D(n1895), .CLK(clk_in), .RSTB(n7254), .Q(
        \FIFO[83][20] ) );
  DFFARX1 \FIFO_reg[83][19]  ( .D(n1894), .CLK(clk_in), .RSTB(n7254), .Q(
        \FIFO[83][19] ) );
  DFFARX1 \FIFO_reg[83][18]  ( .D(n1893), .CLK(clk_in), .RSTB(n7254), .Q(
        \FIFO[83][18] ) );
  DFFARX1 \FIFO_reg[83][17]  ( .D(n1892), .CLK(clk_in), .RSTB(n7255), .Q(
        \FIFO[83][17] ) );
  DFFARX1 \FIFO_reg[83][16]  ( .D(n1891), .CLK(clk_in), .RSTB(n7255), .Q(
        \FIFO[83][16] ) );
  DFFARX1 \FIFO_reg[83][15]  ( .D(n1890), .CLK(clk_in), .RSTB(n7255), .Q(
        \FIFO[83][15] ) );
  DFFARX1 \FIFO_reg[83][14]  ( .D(n1889), .CLK(clk_in), .RSTB(n7255), .Q(
        \FIFO[83][14] ) );
  DFFARX1 \FIFO_reg[83][13]  ( .D(n1888), .CLK(clk_in), .RSTB(n7255), .Q(
        \FIFO[83][13] ) );
  DFFARX1 \FIFO_reg[83][12]  ( .D(n1887), .CLK(clk_in), .RSTB(n7255), .Q(
        \FIFO[83][12] ) );
  DFFARX1 \FIFO_reg[83][11]  ( .D(n1886), .CLK(clk_in), .RSTB(n7255), .Q(
        \FIFO[83][11] ) );
  DFFARX1 \FIFO_reg[83][10]  ( .D(n1885), .CLK(clk_in), .RSTB(n7255), .Q(
        \FIFO[83][10] ) );
  DFFARX1 \FIFO_reg[83][9]  ( .D(n1884), .CLK(clk_in), .RSTB(n7255), .Q(
        \FIFO[83][9] ) );
  DFFARX1 \FIFO_reg[83][8]  ( .D(n1883), .CLK(clk_in), .RSTB(n7255), .Q(
        \FIFO[83][8] ) );
  DFFARX1 \FIFO_reg[83][7]  ( .D(n1882), .CLK(clk_in), .RSTB(n7255), .Q(
        \FIFO[83][7] ) );
  DFFARX1 \FIFO_reg[83][6]  ( .D(n1881), .CLK(clk_in), .RSTB(n7255), .Q(
        \FIFO[83][6] ) );
  DFFARX1 \FIFO_reg[83][5]  ( .D(n1880), .CLK(clk_in), .RSTB(n7255), .Q(
        \FIFO[83][5] ) );
  DFFARX1 \FIFO_reg[83][4]  ( .D(n1879), .CLK(clk_in), .RSTB(n7255), .Q(
        \FIFO[83][4] ) );
  DFFARX1 \FIFO_reg[83][3]  ( .D(n1878), .CLK(clk_in), .RSTB(n7255), .Q(
        \FIFO[83][3] ) );
  DFFARX1 \FIFO_reg[83][2]  ( .D(n1877), .CLK(clk_in), .RSTB(n7255), .Q(
        \FIFO[83][2] ) );
  DFFARX1 \FIFO_reg[83][1]  ( .D(n1876), .CLK(clk_in), .RSTB(n7255), .Q(
        \FIFO[83][1] ) );
  DFFARX1 \FIFO_reg[83][0]  ( .D(n1875), .CLK(clk_in), .RSTB(n7255), .Q(
        \FIFO[83][0] ) );
  DFFARX1 \FIFO_reg[84][31]  ( .D(n1874), .CLK(clk_in), .RSTB(n7256), .Q(
        \FIFO[84][31] ) );
  DFFARX1 \FIFO_reg[84][30]  ( .D(n1873), .CLK(clk_in), .RSTB(n7256), .Q(
        \FIFO[84][30] ) );
  DFFARX1 \FIFO_reg[84][29]  ( .D(n1872), .CLK(clk_in), .RSTB(n7256), .Q(
        \FIFO[84][29] ) );
  DFFARX1 \FIFO_reg[84][28]  ( .D(n1871), .CLK(clk_in), .RSTB(n7256), .Q(
        \FIFO[84][28] ) );
  DFFARX1 \FIFO_reg[84][27]  ( .D(n1870), .CLK(clk_in), .RSTB(n7256), .Q(
        \FIFO[84][27] ) );
  DFFARX1 \FIFO_reg[84][26]  ( .D(n1869), .CLK(clk_in), .RSTB(n7256), .Q(
        \FIFO[84][26] ) );
  DFFARX1 \FIFO_reg[84][25]  ( .D(n1868), .CLK(clk_in), .RSTB(n7256), .Q(
        \FIFO[84][25] ) );
  DFFARX1 \FIFO_reg[84][24]  ( .D(n1867), .CLK(clk_in), .RSTB(n7256), .Q(
        \FIFO[84][24] ) );
  DFFARX1 \FIFO_reg[84][23]  ( .D(n1866), .CLK(clk_in), .RSTB(n7256), .Q(
        \FIFO[84][23] ) );
  DFFARX1 \FIFO_reg[84][22]  ( .D(n1865), .CLK(clk_in), .RSTB(n7256), .Q(
        \FIFO[84][22] ) );
  DFFARX1 \FIFO_reg[84][21]  ( .D(n1864), .CLK(clk_in), .RSTB(n7256), .Q(
        \FIFO[84][21] ) );
  DFFARX1 \FIFO_reg[84][20]  ( .D(n1863), .CLK(clk_in), .RSTB(n7256), .Q(
        \FIFO[84][20] ) );
  DFFARX1 \FIFO_reg[84][19]  ( .D(n1862), .CLK(clk_in), .RSTB(n7256), .Q(
        \FIFO[84][19] ) );
  DFFARX1 \FIFO_reg[84][18]  ( .D(n1861), .CLK(clk_in), .RSTB(n7256), .Q(
        \FIFO[84][18] ) );
  DFFARX1 \FIFO_reg[84][17]  ( .D(n1860), .CLK(clk_in), .RSTB(n7256), .Q(
        \FIFO[84][17] ) );
  DFFARX1 \FIFO_reg[84][16]  ( .D(n1859), .CLK(clk_in), .RSTB(n7256), .Q(
        \FIFO[84][16] ) );
  DFFARX1 \FIFO_reg[84][15]  ( .D(n1858), .CLK(clk_in), .RSTB(n7256), .Q(
        \FIFO[84][15] ) );
  DFFARX1 \FIFO_reg[84][14]  ( .D(n1857), .CLK(clk_in), .RSTB(n7256), .Q(
        \FIFO[84][14] ) );
  DFFARX1 \FIFO_reg[84][13]  ( .D(n1856), .CLK(clk_in), .RSTB(n7257), .Q(
        \FIFO[84][13] ) );
  DFFARX1 \FIFO_reg[84][12]  ( .D(n1855), .CLK(clk_in), .RSTB(n7257), .Q(
        \FIFO[84][12] ) );
  DFFARX1 \FIFO_reg[84][11]  ( .D(n1854), .CLK(clk_in), .RSTB(n7257), .Q(
        \FIFO[84][11] ) );
  DFFARX1 \FIFO_reg[84][10]  ( .D(n1853), .CLK(clk_in), .RSTB(n7257), .Q(
        \FIFO[84][10] ) );
  DFFARX1 \FIFO_reg[84][9]  ( .D(n1852), .CLK(clk_in), .RSTB(n7257), .Q(
        \FIFO[84][9] ) );
  DFFARX1 \FIFO_reg[84][8]  ( .D(n1851), .CLK(clk_in), .RSTB(n7257), .Q(
        \FIFO[84][8] ) );
  DFFARX1 \FIFO_reg[84][7]  ( .D(n1850), .CLK(clk_in), .RSTB(n7257), .Q(
        \FIFO[84][7] ) );
  DFFARX1 \FIFO_reg[84][6]  ( .D(n1849), .CLK(clk_in), .RSTB(n7257), .Q(
        \FIFO[84][6] ) );
  DFFARX1 \FIFO_reg[84][5]  ( .D(n1848), .CLK(clk_in), .RSTB(n7257), .Q(
        \FIFO[84][5] ) );
  DFFARX1 \FIFO_reg[84][4]  ( .D(n1847), .CLK(clk_in), .RSTB(n7257), .Q(
        \FIFO[84][4] ) );
  DFFARX1 \FIFO_reg[84][3]  ( .D(n1846), .CLK(clk_in), .RSTB(n7257), .Q(
        \FIFO[84][3] ) );
  DFFARX1 \FIFO_reg[84][2]  ( .D(n1845), .CLK(clk_in), .RSTB(n7257), .Q(
        \FIFO[84][2] ) );
  DFFARX1 \FIFO_reg[84][1]  ( .D(n1844), .CLK(clk_in), .RSTB(n7257), .Q(
        \FIFO[84][1] ) );
  DFFARX1 \FIFO_reg[84][0]  ( .D(n1843), .CLK(clk_in), .RSTB(n7257), .Q(
        \FIFO[84][0] ) );
  DFFARX1 \FIFO_reg[85][31]  ( .D(n1842), .CLK(clk_in), .RSTB(n7257), .Q(
        \FIFO[85][31] ) );
  DFFARX1 \FIFO_reg[85][30]  ( .D(n1841), .CLK(clk_in), .RSTB(n7257), .Q(
        \FIFO[85][30] ) );
  DFFARX1 \FIFO_reg[85][29]  ( .D(n1840), .CLK(clk_in), .RSTB(n7257), .Q(
        \FIFO[85][29] ) );
  DFFARX1 \FIFO_reg[85][28]  ( .D(n1839), .CLK(clk_in), .RSTB(n7257), .Q(
        \FIFO[85][28] ) );
  DFFARX1 \FIFO_reg[85][27]  ( .D(n1838), .CLK(clk_in), .RSTB(n7258), .Q(
        \FIFO[85][27] ) );
  DFFARX1 \FIFO_reg[85][26]  ( .D(n1837), .CLK(clk_in), .RSTB(n7258), .Q(
        \FIFO[85][26] ) );
  DFFARX1 \FIFO_reg[85][25]  ( .D(n1836), .CLK(clk_in), .RSTB(n7258), .Q(
        \FIFO[85][25] ) );
  DFFARX1 \FIFO_reg[85][24]  ( .D(n1835), .CLK(clk_in), .RSTB(n7258), .Q(
        \FIFO[85][24] ) );
  DFFARX1 \FIFO_reg[85][23]  ( .D(n1834), .CLK(clk_in), .RSTB(n7258), .Q(
        \FIFO[85][23] ) );
  DFFARX1 \FIFO_reg[85][22]  ( .D(n1833), .CLK(clk_in), .RSTB(n7258), .Q(
        \FIFO[85][22] ) );
  DFFARX1 \FIFO_reg[85][21]  ( .D(n1832), .CLK(clk_in), .RSTB(n7258), .Q(
        \FIFO[85][21] ) );
  DFFARX1 \FIFO_reg[85][20]  ( .D(n1831), .CLK(clk_in), .RSTB(n7258), .Q(
        \FIFO[85][20] ) );
  DFFARX1 \FIFO_reg[85][19]  ( .D(n1830), .CLK(clk_in), .RSTB(n7258), .Q(
        \FIFO[85][19] ) );
  DFFARX1 \FIFO_reg[85][18]  ( .D(n1829), .CLK(clk_in), .RSTB(n7258), .Q(
        \FIFO[85][18] ) );
  DFFARX1 \FIFO_reg[85][17]  ( .D(n1828), .CLK(clk_in), .RSTB(n7258), .Q(
        \FIFO[85][17] ) );
  DFFARX1 \FIFO_reg[85][16]  ( .D(n1827), .CLK(clk_in), .RSTB(n7258), .Q(
        \FIFO[85][16] ) );
  DFFARX1 \FIFO_reg[85][15]  ( .D(n1826), .CLK(clk_in), .RSTB(n7258), .Q(
        \FIFO[85][15] ) );
  DFFARX1 \FIFO_reg[85][14]  ( .D(n1825), .CLK(clk_in), .RSTB(n7258), .Q(
        \FIFO[85][14] ) );
  DFFARX1 \FIFO_reg[85][13]  ( .D(n1824), .CLK(clk_in), .RSTB(n7258), .Q(
        \FIFO[85][13] ) );
  DFFARX1 \FIFO_reg[85][12]  ( .D(n1823), .CLK(clk_in), .RSTB(n7258), .Q(
        \FIFO[85][12] ) );
  DFFARX1 \FIFO_reg[85][11]  ( .D(n1822), .CLK(clk_in), .RSTB(n7258), .Q(
        \FIFO[85][11] ) );
  DFFARX1 \FIFO_reg[85][10]  ( .D(n1821), .CLK(clk_in), .RSTB(n7258), .Q(
        \FIFO[85][10] ) );
  DFFARX1 \FIFO_reg[85][9]  ( .D(n1820), .CLK(clk_in), .RSTB(n7259), .Q(
        \FIFO[85][9] ) );
  DFFARX1 \FIFO_reg[85][8]  ( .D(n1819), .CLK(clk_in), .RSTB(n7259), .Q(
        \FIFO[85][8] ) );
  DFFARX1 \FIFO_reg[85][7]  ( .D(n1818), .CLK(clk_in), .RSTB(n7259), .Q(
        \FIFO[85][7] ) );
  DFFARX1 \FIFO_reg[85][6]  ( .D(n1817), .CLK(clk_in), .RSTB(n7259), .Q(
        \FIFO[85][6] ) );
  DFFARX1 \FIFO_reg[85][5]  ( .D(n1816), .CLK(clk_in), .RSTB(n7259), .Q(
        \FIFO[85][5] ) );
  DFFARX1 \FIFO_reg[85][4]  ( .D(n1815), .CLK(clk_in), .RSTB(n7259), .Q(
        \FIFO[85][4] ) );
  DFFARX1 \FIFO_reg[85][3]  ( .D(n1814), .CLK(clk_in), .RSTB(n7259), .Q(
        \FIFO[85][3] ) );
  DFFARX1 \FIFO_reg[85][2]  ( .D(n1813), .CLK(clk_in), .RSTB(n7259), .Q(
        \FIFO[85][2] ) );
  DFFARX1 \FIFO_reg[85][1]  ( .D(n1812), .CLK(clk_in), .RSTB(n7259), .Q(
        \FIFO[85][1] ) );
  DFFARX1 \FIFO_reg[85][0]  ( .D(n1811), .CLK(clk_in), .RSTB(n7259), .Q(
        \FIFO[85][0] ) );
  DFFARX1 \FIFO_reg[86][31]  ( .D(n1810), .CLK(clk_in), .RSTB(n7259), .Q(
        \FIFO[86][31] ) );
  DFFARX1 \FIFO_reg[86][30]  ( .D(n1809), .CLK(clk_in), .RSTB(n7259), .Q(
        \FIFO[86][30] ) );
  DFFARX1 \FIFO_reg[86][29]  ( .D(n1808), .CLK(clk_in), .RSTB(n7259), .Q(
        \FIFO[86][29] ) );
  DFFARX1 \FIFO_reg[86][28]  ( .D(n1807), .CLK(clk_in), .RSTB(n7259), .Q(
        \FIFO[86][28] ) );
  DFFARX1 \FIFO_reg[86][27]  ( .D(n1806), .CLK(clk_in), .RSTB(n7259), .Q(
        \FIFO[86][27] ) );
  DFFARX1 \FIFO_reg[86][26]  ( .D(n1805), .CLK(clk_in), .RSTB(n7259), .Q(
        \FIFO[86][26] ) );
  DFFARX1 \FIFO_reg[86][25]  ( .D(n1804), .CLK(clk_in), .RSTB(n7259), .Q(
        \FIFO[86][25] ) );
  DFFARX1 \FIFO_reg[86][24]  ( .D(n1803), .CLK(clk_in), .RSTB(n7259), .Q(
        \FIFO[86][24] ) );
  DFFARX1 \FIFO_reg[86][23]  ( .D(n1802), .CLK(clk_in), .RSTB(n7260), .Q(
        \FIFO[86][23] ) );
  DFFARX1 \FIFO_reg[86][22]  ( .D(n1801), .CLK(clk_in), .RSTB(n7260), .Q(
        \FIFO[86][22] ) );
  DFFARX1 \FIFO_reg[86][21]  ( .D(n1800), .CLK(clk_in), .RSTB(n7260), .Q(
        \FIFO[86][21] ) );
  DFFARX1 \FIFO_reg[86][20]  ( .D(n1799), .CLK(clk_in), .RSTB(n7260), .Q(
        \FIFO[86][20] ) );
  DFFARX1 \FIFO_reg[86][19]  ( .D(n1798), .CLK(clk_in), .RSTB(n7260), .Q(
        \FIFO[86][19] ) );
  DFFARX1 \FIFO_reg[86][18]  ( .D(n1797), .CLK(clk_in), .RSTB(n7260), .Q(
        \FIFO[86][18] ) );
  DFFARX1 \FIFO_reg[86][17]  ( .D(n1796), .CLK(clk_in), .RSTB(n7260), .Q(
        \FIFO[86][17] ) );
  DFFARX1 \FIFO_reg[86][16]  ( .D(n1795), .CLK(clk_in), .RSTB(n7260), .Q(
        \FIFO[86][16] ) );
  DFFARX1 \FIFO_reg[86][15]  ( .D(n1794), .CLK(clk_in), .RSTB(n7260), .Q(
        \FIFO[86][15] ) );
  DFFARX1 \FIFO_reg[86][14]  ( .D(n1793), .CLK(clk_in), .RSTB(n7260), .Q(
        \FIFO[86][14] ) );
  DFFARX1 \FIFO_reg[86][13]  ( .D(n1792), .CLK(clk_in), .RSTB(n7260), .Q(
        \FIFO[86][13] ) );
  DFFARX1 \FIFO_reg[86][12]  ( .D(n1791), .CLK(clk_in), .RSTB(n7260), .Q(
        \FIFO[86][12] ) );
  DFFARX1 \FIFO_reg[86][11]  ( .D(n1790), .CLK(clk_in), .RSTB(n7260), .Q(
        \FIFO[86][11] ) );
  DFFARX1 \FIFO_reg[86][10]  ( .D(n1789), .CLK(clk_in), .RSTB(n7260), .Q(
        \FIFO[86][10] ) );
  DFFARX1 \FIFO_reg[86][9]  ( .D(n1788), .CLK(clk_in), .RSTB(n7260), .Q(
        \FIFO[86][9] ) );
  DFFARX1 \FIFO_reg[86][8]  ( .D(n1787), .CLK(clk_in), .RSTB(n7260), .Q(
        \FIFO[86][8] ) );
  DFFARX1 \FIFO_reg[86][7]  ( .D(n1786), .CLK(clk_in), .RSTB(n7260), .Q(
        \FIFO[86][7] ) );
  DFFARX1 \FIFO_reg[86][6]  ( .D(n1785), .CLK(clk_in), .RSTB(n7260), .Q(
        \FIFO[86][6] ) );
  DFFARX1 \FIFO_reg[86][5]  ( .D(n1784), .CLK(clk_in), .RSTB(n7261), .Q(
        \FIFO[86][5] ) );
  DFFARX1 \FIFO_reg[86][4]  ( .D(n1783), .CLK(clk_in), .RSTB(n7261), .Q(
        \FIFO[86][4] ) );
  DFFARX1 \FIFO_reg[86][3]  ( .D(n1782), .CLK(clk_in), .RSTB(n7261), .Q(
        \FIFO[86][3] ) );
  DFFARX1 \FIFO_reg[86][2]  ( .D(n1781), .CLK(clk_in), .RSTB(n7261), .Q(
        \FIFO[86][2] ) );
  DFFARX1 \FIFO_reg[86][1]  ( .D(n1780), .CLK(clk_in), .RSTB(n7261), .Q(
        \FIFO[86][1] ) );
  DFFARX1 \FIFO_reg[86][0]  ( .D(n1779), .CLK(clk_in), .RSTB(n7261), .Q(
        \FIFO[86][0] ) );
  DFFARX1 \FIFO_reg[87][31]  ( .D(n1778), .CLK(clk_in), .RSTB(n7261), .Q(
        \FIFO[87][31] ) );
  DFFARX1 \FIFO_reg[87][30]  ( .D(n1777), .CLK(clk_in), .RSTB(n7261), .Q(
        \FIFO[87][30] ) );
  DFFARX1 \FIFO_reg[87][29]  ( .D(n1776), .CLK(clk_in), .RSTB(n7261), .Q(
        \FIFO[87][29] ) );
  DFFARX1 \FIFO_reg[87][28]  ( .D(n1775), .CLK(clk_in), .RSTB(n7261), .Q(
        \FIFO[87][28] ) );
  DFFARX1 \FIFO_reg[87][27]  ( .D(n1774), .CLK(clk_in), .RSTB(n7261), .Q(
        \FIFO[87][27] ) );
  DFFARX1 \FIFO_reg[87][26]  ( .D(n1773), .CLK(clk_in), .RSTB(n7261), .Q(
        \FIFO[87][26] ) );
  DFFARX1 \FIFO_reg[87][25]  ( .D(n1772), .CLK(clk_in), .RSTB(n7261), .Q(
        \FIFO[87][25] ) );
  DFFARX1 \FIFO_reg[87][24]  ( .D(n1771), .CLK(clk_in), .RSTB(n7261), .Q(
        \FIFO[87][24] ) );
  DFFARX1 \FIFO_reg[87][23]  ( .D(n1770), .CLK(clk_in), .RSTB(n7261), .Q(
        \FIFO[87][23] ) );
  DFFARX1 \FIFO_reg[87][22]  ( .D(n1769), .CLK(clk_in), .RSTB(n7261), .Q(
        \FIFO[87][22] ) );
  DFFARX1 \FIFO_reg[87][21]  ( .D(n1768), .CLK(clk_in), .RSTB(n7261), .Q(
        \FIFO[87][21] ) );
  DFFARX1 \FIFO_reg[87][20]  ( .D(n1767), .CLK(clk_in), .RSTB(n7261), .Q(
        \FIFO[87][20] ) );
  DFFARX1 \FIFO_reg[87][19]  ( .D(n1766), .CLK(clk_in), .RSTB(n7262), .Q(
        \FIFO[87][19] ) );
  DFFARX1 \FIFO_reg[87][18]  ( .D(n1765), .CLK(clk_in), .RSTB(n7262), .Q(
        \FIFO[87][18] ) );
  DFFARX1 \FIFO_reg[87][17]  ( .D(n1764), .CLK(clk_in), .RSTB(n7262), .Q(
        \FIFO[87][17] ) );
  DFFARX1 \FIFO_reg[87][16]  ( .D(n1763), .CLK(clk_in), .RSTB(n7262), .Q(
        \FIFO[87][16] ) );
  DFFARX1 \FIFO_reg[87][15]  ( .D(n1762), .CLK(clk_in), .RSTB(n7262), .Q(
        \FIFO[87][15] ) );
  DFFARX1 \FIFO_reg[87][14]  ( .D(n1761), .CLK(clk_in), .RSTB(n7262), .Q(
        \FIFO[87][14] ) );
  DFFARX1 \FIFO_reg[87][13]  ( .D(n1760), .CLK(clk_in), .RSTB(n7262), .Q(
        \FIFO[87][13] ) );
  DFFARX1 \FIFO_reg[87][12]  ( .D(n1759), .CLK(clk_in), .RSTB(n7262), .Q(
        \FIFO[87][12] ) );
  DFFARX1 \FIFO_reg[87][11]  ( .D(n1758), .CLK(clk_in), .RSTB(n7262), .Q(
        \FIFO[87][11] ) );
  DFFARX1 \FIFO_reg[87][10]  ( .D(n1757), .CLK(clk_in), .RSTB(n7262), .Q(
        \FIFO[87][10] ) );
  DFFARX1 \FIFO_reg[87][9]  ( .D(n1756), .CLK(clk_in), .RSTB(n7262), .Q(
        \FIFO[87][9] ) );
  DFFARX1 \FIFO_reg[87][8]  ( .D(n1755), .CLK(clk_in), .RSTB(n7262), .Q(
        \FIFO[87][8] ) );
  DFFARX1 \FIFO_reg[87][7]  ( .D(n1754), .CLK(clk_in), .RSTB(n7262), .Q(
        \FIFO[87][7] ) );
  DFFARX1 \FIFO_reg[87][6]  ( .D(n1753), .CLK(clk_in), .RSTB(n7262), .Q(
        \FIFO[87][6] ) );
  DFFARX1 \FIFO_reg[87][5]  ( .D(n1752), .CLK(clk_in), .RSTB(n7262), .Q(
        \FIFO[87][5] ) );
  DFFARX1 \FIFO_reg[87][4]  ( .D(n1751), .CLK(clk_in), .RSTB(n7262), .Q(
        \FIFO[87][4] ) );
  DFFARX1 \FIFO_reg[87][3]  ( .D(n1750), .CLK(clk_in), .RSTB(n7262), .Q(
        \FIFO[87][3] ) );
  DFFARX1 \FIFO_reg[87][2]  ( .D(n1749), .CLK(clk_in), .RSTB(n7262), .Q(
        \FIFO[87][2] ) );
  DFFARX1 \FIFO_reg[87][1]  ( .D(n1748), .CLK(clk_in), .RSTB(n7263), .Q(
        \FIFO[87][1] ) );
  DFFARX1 \FIFO_reg[87][0]  ( .D(n1747), .CLK(clk_in), .RSTB(n7263), .Q(
        \FIFO[87][0] ) );
  DFFARX1 \FIFO_reg[88][31]  ( .D(n1746), .CLK(clk_in), .RSTB(n7263), .Q(
        \FIFO[88][31] ) );
  DFFARX1 \FIFO_reg[88][30]  ( .D(n1745), .CLK(clk_in), .RSTB(n7263), .Q(
        \FIFO[88][30] ) );
  DFFARX1 \FIFO_reg[88][29]  ( .D(n1744), .CLK(clk_in), .RSTB(n7263), .Q(
        \FIFO[88][29] ) );
  DFFARX1 \FIFO_reg[88][28]  ( .D(n1743), .CLK(clk_in), .RSTB(n7263), .Q(
        \FIFO[88][28] ) );
  DFFARX1 \FIFO_reg[88][27]  ( .D(n1742), .CLK(clk_in), .RSTB(n7263), .Q(
        \FIFO[88][27] ) );
  DFFARX1 \FIFO_reg[88][26]  ( .D(n1741), .CLK(clk_in), .RSTB(n7263), .Q(
        \FIFO[88][26] ) );
  DFFARX1 \FIFO_reg[88][25]  ( .D(n1740), .CLK(clk_in), .RSTB(n7263), .Q(
        \FIFO[88][25] ) );
  DFFARX1 \FIFO_reg[88][24]  ( .D(n1739), .CLK(clk_in), .RSTB(n7263), .Q(
        \FIFO[88][24] ) );
  DFFARX1 \FIFO_reg[88][23]  ( .D(n1738), .CLK(clk_in), .RSTB(n7263), .Q(
        \FIFO[88][23] ) );
  DFFARX1 \FIFO_reg[88][22]  ( .D(n1737), .CLK(clk_in), .RSTB(n7263), .Q(
        \FIFO[88][22] ) );
  DFFARX1 \FIFO_reg[88][21]  ( .D(n1736), .CLK(clk_in), .RSTB(n7263), .Q(
        \FIFO[88][21] ) );
  DFFARX1 \FIFO_reg[88][20]  ( .D(n1735), .CLK(clk_in), .RSTB(n7263), .Q(
        \FIFO[88][20] ) );
  DFFARX1 \FIFO_reg[88][19]  ( .D(n1734), .CLK(clk_in), .RSTB(n7263), .Q(
        \FIFO[88][19] ) );
  DFFARX1 \FIFO_reg[88][18]  ( .D(n1733), .CLK(clk_in), .RSTB(n7263), .Q(
        \FIFO[88][18] ) );
  DFFARX1 \FIFO_reg[88][17]  ( .D(n1732), .CLK(clk_in), .RSTB(n7263), .Q(
        \FIFO[88][17] ) );
  DFFARX1 \FIFO_reg[88][16]  ( .D(n1731), .CLK(clk_in), .RSTB(n7263), .Q(
        \FIFO[88][16] ) );
  DFFARX1 \FIFO_reg[88][15]  ( .D(n1730), .CLK(clk_in), .RSTB(n7264), .Q(
        \FIFO[88][15] ) );
  DFFARX1 \FIFO_reg[88][14]  ( .D(n1729), .CLK(clk_in), .RSTB(n7264), .Q(
        \FIFO[88][14] ) );
  DFFARX1 \FIFO_reg[88][13]  ( .D(n1728), .CLK(clk_in), .RSTB(n7264), .Q(
        \FIFO[88][13] ) );
  DFFARX1 \FIFO_reg[88][12]  ( .D(n1727), .CLK(clk_in), .RSTB(n7264), .Q(
        \FIFO[88][12] ) );
  DFFARX1 \FIFO_reg[88][11]  ( .D(n1726), .CLK(clk_in), .RSTB(n7264), .Q(
        \FIFO[88][11] ) );
  DFFARX1 \FIFO_reg[88][10]  ( .D(n1725), .CLK(clk_in), .RSTB(n7264), .Q(
        \FIFO[88][10] ) );
  DFFARX1 \FIFO_reg[88][9]  ( .D(n1724), .CLK(clk_in), .RSTB(n7264), .Q(
        \FIFO[88][9] ) );
  DFFARX1 \FIFO_reg[88][8]  ( .D(n1723), .CLK(clk_in), .RSTB(n7264), .Q(
        \FIFO[88][8] ) );
  DFFARX1 \FIFO_reg[88][7]  ( .D(n1722), .CLK(clk_in), .RSTB(n7264), .Q(
        \FIFO[88][7] ) );
  DFFARX1 \FIFO_reg[88][6]  ( .D(n1721), .CLK(clk_in), .RSTB(n7264), .Q(
        \FIFO[88][6] ) );
  DFFARX1 \FIFO_reg[88][5]  ( .D(n1720), .CLK(clk_in), .RSTB(n7264), .Q(
        \FIFO[88][5] ) );
  DFFARX1 \FIFO_reg[88][4]  ( .D(n1719), .CLK(clk_in), .RSTB(n7264), .Q(
        \FIFO[88][4] ) );
  DFFARX1 \FIFO_reg[88][3]  ( .D(n1718), .CLK(clk_in), .RSTB(n7264), .Q(
        \FIFO[88][3] ) );
  DFFARX1 \FIFO_reg[88][2]  ( .D(n1717), .CLK(clk_in), .RSTB(n7264), .Q(
        \FIFO[88][2] ) );
  DFFARX1 \FIFO_reg[88][1]  ( .D(n1716), .CLK(clk_in), .RSTB(n7264), .Q(
        \FIFO[88][1] ) );
  DFFARX1 \FIFO_reg[88][0]  ( .D(n1715), .CLK(clk_in), .RSTB(n7264), .Q(
        \FIFO[88][0] ) );
  DFFARX1 \FIFO_reg[89][31]  ( .D(n1714), .CLK(clk_in), .RSTB(n7264), .Q(
        \FIFO[89][31] ) );
  DFFARX1 \FIFO_reg[89][30]  ( .D(n1713), .CLK(clk_in), .RSTB(n7264), .Q(
        \FIFO[89][30] ) );
  DFFARX1 \FIFO_reg[89][29]  ( .D(n1712), .CLK(clk_in), .RSTB(n7265), .Q(
        \FIFO[89][29] ) );
  DFFARX1 \FIFO_reg[89][28]  ( .D(n1711), .CLK(clk_in), .RSTB(n7265), .Q(
        \FIFO[89][28] ) );
  DFFARX1 \FIFO_reg[89][27]  ( .D(n1710), .CLK(clk_in), .RSTB(n7265), .Q(
        \FIFO[89][27] ) );
  DFFARX1 \FIFO_reg[89][26]  ( .D(n1709), .CLK(clk_in), .RSTB(n7265), .Q(
        \FIFO[89][26] ) );
  DFFARX1 \FIFO_reg[89][25]  ( .D(n1708), .CLK(clk_in), .RSTB(n7265), .Q(
        \FIFO[89][25] ) );
  DFFARX1 \FIFO_reg[89][24]  ( .D(n1707), .CLK(clk_in), .RSTB(n7265), .Q(
        \FIFO[89][24] ) );
  DFFARX1 \FIFO_reg[89][23]  ( .D(n1706), .CLK(clk_in), .RSTB(n7265), .Q(
        \FIFO[89][23] ) );
  DFFARX1 \FIFO_reg[89][22]  ( .D(n1705), .CLK(clk_in), .RSTB(n7265), .Q(
        \FIFO[89][22] ) );
  DFFARX1 \FIFO_reg[89][21]  ( .D(n1704), .CLK(clk_in), .RSTB(n7265), .Q(
        \FIFO[89][21] ) );
  DFFARX1 \FIFO_reg[89][20]  ( .D(n1703), .CLK(clk_in), .RSTB(n7265), .Q(
        \FIFO[89][20] ) );
  DFFARX1 \FIFO_reg[89][19]  ( .D(n1702), .CLK(clk_in), .RSTB(n7265), .Q(
        \FIFO[89][19] ) );
  DFFARX1 \FIFO_reg[89][18]  ( .D(n1701), .CLK(clk_in), .RSTB(n7265), .Q(
        \FIFO[89][18] ) );
  DFFARX1 \FIFO_reg[89][17]  ( .D(n1700), .CLK(clk_in), .RSTB(n7265), .Q(
        \FIFO[89][17] ) );
  DFFARX1 \FIFO_reg[89][16]  ( .D(n1699), .CLK(clk_in), .RSTB(n7265), .Q(
        \FIFO[89][16] ) );
  DFFARX1 \FIFO_reg[89][15]  ( .D(n1698), .CLK(clk_in), .RSTB(n7265), .Q(
        \FIFO[89][15] ) );
  DFFARX1 \FIFO_reg[89][14]  ( .D(n1697), .CLK(clk_in), .RSTB(n7265), .Q(
        \FIFO[89][14] ) );
  DFFARX1 \FIFO_reg[89][13]  ( .D(n1696), .CLK(clk_in), .RSTB(n7265), .Q(
        \FIFO[89][13] ) );
  DFFARX1 \FIFO_reg[89][12]  ( .D(n1695), .CLK(clk_in), .RSTB(n7265), .Q(
        \FIFO[89][12] ) );
  DFFARX1 \FIFO_reg[89][11]  ( .D(n1694), .CLK(clk_in), .RSTB(n7266), .Q(
        \FIFO[89][11] ) );
  DFFARX1 \FIFO_reg[89][10]  ( .D(n1693), .CLK(clk_in), .RSTB(n7266), .Q(
        \FIFO[89][10] ) );
  DFFARX1 \FIFO_reg[89][9]  ( .D(n1692), .CLK(clk_in), .RSTB(n7266), .Q(
        \FIFO[89][9] ) );
  DFFARX1 \FIFO_reg[89][8]  ( .D(n1691), .CLK(clk_in), .RSTB(n7266), .Q(
        \FIFO[89][8] ) );
  DFFARX1 \FIFO_reg[89][7]  ( .D(n1690), .CLK(clk_in), .RSTB(n7266), .Q(
        \FIFO[89][7] ) );
  DFFARX1 \FIFO_reg[89][6]  ( .D(n1689), .CLK(clk_in), .RSTB(n7266), .Q(
        \FIFO[89][6] ) );
  DFFARX1 \FIFO_reg[89][5]  ( .D(n1688), .CLK(clk_in), .RSTB(n7266), .Q(
        \FIFO[89][5] ) );
  DFFARX1 \FIFO_reg[89][4]  ( .D(n1687), .CLK(clk_in), .RSTB(n7266), .Q(
        \FIFO[89][4] ) );
  DFFARX1 \FIFO_reg[89][3]  ( .D(n1686), .CLK(clk_in), .RSTB(n7266), .Q(
        \FIFO[89][3] ) );
  DFFARX1 \FIFO_reg[89][2]  ( .D(n1685), .CLK(clk_in), .RSTB(n7266), .Q(
        \FIFO[89][2] ) );
  DFFARX1 \FIFO_reg[89][1]  ( .D(n1684), .CLK(clk_in), .RSTB(n7266), .Q(
        \FIFO[89][1] ) );
  DFFARX1 \FIFO_reg[89][0]  ( .D(n1683), .CLK(clk_in), .RSTB(n7266), .Q(
        \FIFO[89][0] ) );
  DFFARX1 \FIFO_reg[90][31]  ( .D(n1682), .CLK(clk_in), .RSTB(n7266), .Q(
        \FIFO[90][31] ) );
  DFFARX1 \FIFO_reg[90][30]  ( .D(n1681), .CLK(clk_in), .RSTB(n7266), .Q(
        \FIFO[90][30] ) );
  DFFARX1 \FIFO_reg[90][29]  ( .D(n1680), .CLK(clk_in), .RSTB(n7266), .Q(
        \FIFO[90][29] ) );
  DFFARX1 \FIFO_reg[90][28]  ( .D(n1679), .CLK(clk_in), .RSTB(n7266), .Q(
        \FIFO[90][28] ) );
  DFFARX1 \FIFO_reg[90][27]  ( .D(n1678), .CLK(clk_in), .RSTB(n7266), .Q(
        \FIFO[90][27] ) );
  DFFARX1 \FIFO_reg[90][26]  ( .D(n1677), .CLK(clk_in), .RSTB(n7266), .Q(
        \FIFO[90][26] ) );
  DFFARX1 \FIFO_reg[90][25]  ( .D(n1676), .CLK(clk_in), .RSTB(n7267), .Q(
        \FIFO[90][25] ) );
  DFFARX1 \FIFO_reg[90][24]  ( .D(n1675), .CLK(clk_in), .RSTB(n7267), .Q(
        \FIFO[90][24] ) );
  DFFARX1 \FIFO_reg[90][23]  ( .D(n1674), .CLK(clk_in), .RSTB(n7267), .Q(
        \FIFO[90][23] ) );
  DFFARX1 \FIFO_reg[90][22]  ( .D(n1673), .CLK(clk_in), .RSTB(n7267), .Q(
        \FIFO[90][22] ) );
  DFFARX1 \FIFO_reg[90][21]  ( .D(n1672), .CLK(clk_in), .RSTB(n7267), .Q(
        \FIFO[90][21] ) );
  DFFARX1 \FIFO_reg[90][20]  ( .D(n1671), .CLK(clk_in), .RSTB(n7267), .Q(
        \FIFO[90][20] ) );
  DFFARX1 \FIFO_reg[90][19]  ( .D(n1670), .CLK(clk_in), .RSTB(n7267), .Q(
        \FIFO[90][19] ) );
  DFFARX1 \FIFO_reg[90][18]  ( .D(n1669), .CLK(clk_in), .RSTB(n7267), .Q(
        \FIFO[90][18] ) );
  DFFARX1 \FIFO_reg[90][17]  ( .D(n1668), .CLK(clk_in), .RSTB(n7267), .Q(
        \FIFO[90][17] ) );
  DFFARX1 \FIFO_reg[90][16]  ( .D(n1667), .CLK(clk_in), .RSTB(n7267), .Q(
        \FIFO[90][16] ) );
  DFFARX1 \FIFO_reg[90][15]  ( .D(n1666), .CLK(clk_in), .RSTB(n7267), .Q(
        \FIFO[90][15] ) );
  DFFARX1 \FIFO_reg[90][14]  ( .D(n1665), .CLK(clk_in), .RSTB(n7267), .Q(
        \FIFO[90][14] ) );
  DFFARX1 \FIFO_reg[90][13]  ( .D(n1664), .CLK(clk_in), .RSTB(n7267), .Q(
        \FIFO[90][13] ) );
  DFFARX1 \FIFO_reg[90][12]  ( .D(n1663), .CLK(clk_in), .RSTB(n7267), .Q(
        \FIFO[90][12] ) );
  DFFARX1 \FIFO_reg[90][11]  ( .D(n1662), .CLK(clk_in), .RSTB(n7267), .Q(
        \FIFO[90][11] ) );
  DFFARX1 \FIFO_reg[90][10]  ( .D(n1661), .CLK(clk_in), .RSTB(n7267), .Q(
        \FIFO[90][10] ) );
  DFFARX1 \FIFO_reg[90][9]  ( .D(n1660), .CLK(clk_in), .RSTB(n7267), .Q(
        \FIFO[90][9] ) );
  DFFARX1 \FIFO_reg[90][8]  ( .D(n1659), .CLK(clk_in), .RSTB(n7267), .Q(
        \FIFO[90][8] ) );
  DFFARX1 \FIFO_reg[90][7]  ( .D(n1658), .CLK(clk_in), .RSTB(n7268), .Q(
        \FIFO[90][7] ) );
  DFFARX1 \FIFO_reg[90][6]  ( .D(n1657), .CLK(clk_in), .RSTB(n7268), .Q(
        \FIFO[90][6] ) );
  DFFARX1 \FIFO_reg[90][5]  ( .D(n1656), .CLK(clk_in), .RSTB(n7268), .Q(
        \FIFO[90][5] ) );
  DFFARX1 \FIFO_reg[90][4]  ( .D(n1655), .CLK(clk_in), .RSTB(n7268), .Q(
        \FIFO[90][4] ) );
  DFFARX1 \FIFO_reg[90][3]  ( .D(n1654), .CLK(clk_in), .RSTB(n7268), .Q(
        \FIFO[90][3] ) );
  DFFARX1 \FIFO_reg[90][2]  ( .D(n1653), .CLK(clk_in), .RSTB(n7268), .Q(
        \FIFO[90][2] ) );
  DFFARX1 \FIFO_reg[90][1]  ( .D(n1652), .CLK(clk_in), .RSTB(n7268), .Q(
        \FIFO[90][1] ) );
  DFFARX1 \FIFO_reg[90][0]  ( .D(n1651), .CLK(clk_in), .RSTB(n7268), .Q(
        \FIFO[90][0] ) );
  DFFARX1 \FIFO_reg[91][31]  ( .D(n1650), .CLK(clk_in), .RSTB(n7268), .Q(
        \FIFO[91][31] ) );
  DFFARX1 \FIFO_reg[91][30]  ( .D(n1649), .CLK(clk_in), .RSTB(n7268), .Q(
        \FIFO[91][30] ) );
  DFFARX1 \FIFO_reg[91][29]  ( .D(n1648), .CLK(clk_in), .RSTB(n7268), .Q(
        \FIFO[91][29] ) );
  DFFARX1 \FIFO_reg[91][28]  ( .D(n1647), .CLK(clk_in), .RSTB(n7268), .Q(
        \FIFO[91][28] ) );
  DFFARX1 \FIFO_reg[91][27]  ( .D(n1646), .CLK(clk_in), .RSTB(n7268), .Q(
        \FIFO[91][27] ) );
  DFFARX1 \FIFO_reg[91][26]  ( .D(n1645), .CLK(clk_in), .RSTB(n7268), .Q(
        \FIFO[91][26] ) );
  DFFARX1 \FIFO_reg[91][25]  ( .D(n1644), .CLK(clk_in), .RSTB(n7268), .Q(
        \FIFO[91][25] ) );
  DFFARX1 \FIFO_reg[91][24]  ( .D(n1643), .CLK(clk_in), .RSTB(n7268), .Q(
        \FIFO[91][24] ) );
  DFFARX1 \FIFO_reg[91][23]  ( .D(n1642), .CLK(clk_in), .RSTB(n7268), .Q(
        \FIFO[91][23] ) );
  DFFARX1 \FIFO_reg[91][22]  ( .D(n1641), .CLK(clk_in), .RSTB(n7268), .Q(
        \FIFO[91][22] ) );
  DFFARX1 \FIFO_reg[91][21]  ( .D(n1640), .CLK(clk_in), .RSTB(n7269), .Q(
        \FIFO[91][21] ) );
  DFFARX1 \FIFO_reg[91][20]  ( .D(n1639), .CLK(clk_in), .RSTB(n7269), .Q(
        \FIFO[91][20] ) );
  DFFARX1 \FIFO_reg[91][19]  ( .D(n1638), .CLK(clk_in), .RSTB(n7269), .Q(
        \FIFO[91][19] ) );
  DFFARX1 \FIFO_reg[91][18]  ( .D(n1637), .CLK(clk_in), .RSTB(n7269), .Q(
        \FIFO[91][18] ) );
  DFFARX1 \FIFO_reg[91][17]  ( .D(n1636), .CLK(clk_in), .RSTB(n7269), .Q(
        \FIFO[91][17] ) );
  DFFARX1 \FIFO_reg[91][16]  ( .D(n1635), .CLK(clk_in), .RSTB(n7269), .Q(
        \FIFO[91][16] ) );
  DFFARX1 \FIFO_reg[91][15]  ( .D(n1634), .CLK(clk_in), .RSTB(n7269), .Q(
        \FIFO[91][15] ) );
  DFFARX1 \FIFO_reg[91][14]  ( .D(n1633), .CLK(clk_in), .RSTB(n7269), .Q(
        \FIFO[91][14] ) );
  DFFARX1 \FIFO_reg[91][13]  ( .D(n1632), .CLK(clk_in), .RSTB(n7269), .Q(
        \FIFO[91][13] ) );
  DFFARX1 \FIFO_reg[91][12]  ( .D(n1631), .CLK(clk_in), .RSTB(n7269), .Q(
        \FIFO[91][12] ) );
  DFFARX1 \FIFO_reg[91][11]  ( .D(n1630), .CLK(clk_in), .RSTB(n7269), .Q(
        \FIFO[91][11] ) );
  DFFARX1 \FIFO_reg[91][10]  ( .D(n1629), .CLK(clk_in), .RSTB(n7269), .Q(
        \FIFO[91][10] ) );
  DFFARX1 \FIFO_reg[91][9]  ( .D(n1628), .CLK(clk_in), .RSTB(n7269), .Q(
        \FIFO[91][9] ) );
  DFFARX1 \FIFO_reg[91][8]  ( .D(n1627), .CLK(clk_in), .RSTB(n7269), .Q(
        \FIFO[91][8] ) );
  DFFARX1 \FIFO_reg[91][7]  ( .D(n1626), .CLK(clk_in), .RSTB(n7269), .Q(
        \FIFO[91][7] ) );
  DFFARX1 \FIFO_reg[91][6]  ( .D(n1625), .CLK(clk_in), .RSTB(n7269), .Q(
        \FIFO[91][6] ) );
  DFFARX1 \FIFO_reg[91][5]  ( .D(n1624), .CLK(clk_in), .RSTB(n7269), .Q(
        \FIFO[91][5] ) );
  DFFARX1 \FIFO_reg[91][4]  ( .D(n1623), .CLK(clk_in), .RSTB(n7269), .Q(
        \FIFO[91][4] ) );
  DFFARX1 \FIFO_reg[91][3]  ( .D(n1622), .CLK(clk_in), .RSTB(n7270), .Q(
        \FIFO[91][3] ) );
  DFFARX1 \FIFO_reg[91][2]  ( .D(n1621), .CLK(clk_in), .RSTB(n7270), .Q(
        \FIFO[91][2] ) );
  DFFARX1 \FIFO_reg[91][1]  ( .D(n1620), .CLK(clk_in), .RSTB(n7270), .Q(
        \FIFO[91][1] ) );
  DFFARX1 \FIFO_reg[91][0]  ( .D(n1619), .CLK(clk_in), .RSTB(n7270), .Q(
        \FIFO[91][0] ) );
  DFFARX1 \FIFO_reg[92][31]  ( .D(n1618), .CLK(clk_in), .RSTB(n7270), .Q(
        \FIFO[92][31] ) );
  DFFARX1 \FIFO_reg[92][30]  ( .D(n1617), .CLK(clk_in), .RSTB(n7270), .Q(
        \FIFO[92][30] ) );
  DFFARX1 \FIFO_reg[92][29]  ( .D(n1616), .CLK(clk_in), .RSTB(n7270), .Q(
        \FIFO[92][29] ) );
  DFFARX1 \FIFO_reg[92][28]  ( .D(n1615), .CLK(clk_in), .RSTB(n7270), .Q(
        \FIFO[92][28] ) );
  DFFARX1 \FIFO_reg[92][27]  ( .D(n1614), .CLK(clk_in), .RSTB(n7270), .Q(
        \FIFO[92][27] ) );
  DFFARX1 \FIFO_reg[92][26]  ( .D(n1613), .CLK(clk_in), .RSTB(n7270), .Q(
        \FIFO[92][26] ) );
  DFFARX1 \FIFO_reg[92][25]  ( .D(n1612), .CLK(clk_in), .RSTB(n7270), .Q(
        \FIFO[92][25] ) );
  DFFARX1 \FIFO_reg[92][24]  ( .D(n1611), .CLK(clk_in), .RSTB(n7270), .Q(
        \FIFO[92][24] ) );
  DFFARX1 \FIFO_reg[92][23]  ( .D(n1610), .CLK(clk_in), .RSTB(n7270), .Q(
        \FIFO[92][23] ) );
  DFFARX1 \FIFO_reg[92][22]  ( .D(n1609), .CLK(clk_in), .RSTB(n7270), .Q(
        \FIFO[92][22] ) );
  DFFARX1 \FIFO_reg[92][21]  ( .D(n1608), .CLK(clk_in), .RSTB(n7270), .Q(
        \FIFO[92][21] ) );
  DFFARX1 \FIFO_reg[92][20]  ( .D(n1607), .CLK(clk_in), .RSTB(n7270), .Q(
        \FIFO[92][20] ) );
  DFFARX1 \FIFO_reg[92][19]  ( .D(n1606), .CLK(clk_in), .RSTB(n7270), .Q(
        \FIFO[92][19] ) );
  DFFARX1 \FIFO_reg[92][18]  ( .D(n1605), .CLK(clk_in), .RSTB(n7270), .Q(
        \FIFO[92][18] ) );
  DFFARX1 \FIFO_reg[92][17]  ( .D(n1604), .CLK(clk_in), .RSTB(n7271), .Q(
        \FIFO[92][17] ) );
  DFFARX1 \FIFO_reg[92][16]  ( .D(n1603), .CLK(clk_in), .RSTB(n7271), .Q(
        \FIFO[92][16] ) );
  DFFARX1 \FIFO_reg[92][15]  ( .D(n1602), .CLK(clk_in), .RSTB(n7271), .Q(
        \FIFO[92][15] ) );
  DFFARX1 \FIFO_reg[92][14]  ( .D(n1601), .CLK(clk_in), .RSTB(n7271), .Q(
        \FIFO[92][14] ) );
  DFFARX1 \FIFO_reg[92][13]  ( .D(n1600), .CLK(clk_in), .RSTB(n7271), .Q(
        \FIFO[92][13] ) );
  DFFARX1 \FIFO_reg[92][12]  ( .D(n1599), .CLK(clk_in), .RSTB(n7271), .Q(
        \FIFO[92][12] ) );
  DFFARX1 \FIFO_reg[92][11]  ( .D(n1598), .CLK(clk_in), .RSTB(n7271), .Q(
        \FIFO[92][11] ) );
  DFFARX1 \FIFO_reg[92][10]  ( .D(n1597), .CLK(clk_in), .RSTB(n7271), .Q(
        \FIFO[92][10] ) );
  DFFARX1 \FIFO_reg[92][9]  ( .D(n1596), .CLK(clk_in), .RSTB(n7271), .Q(
        \FIFO[92][9] ) );
  DFFARX1 \FIFO_reg[92][8]  ( .D(n1595), .CLK(clk_in), .RSTB(n7271), .Q(
        \FIFO[92][8] ) );
  DFFARX1 \FIFO_reg[92][7]  ( .D(n1594), .CLK(clk_in), .RSTB(n7271), .Q(
        \FIFO[92][7] ) );
  DFFARX1 \FIFO_reg[92][6]  ( .D(n1593), .CLK(clk_in), .RSTB(n7271), .Q(
        \FIFO[92][6] ) );
  DFFARX1 \FIFO_reg[92][5]  ( .D(n1592), .CLK(clk_in), .RSTB(n7271), .Q(
        \FIFO[92][5] ) );
  DFFARX1 \FIFO_reg[92][4]  ( .D(n1591), .CLK(clk_in), .RSTB(n7271), .Q(
        \FIFO[92][4] ) );
  DFFARX1 \FIFO_reg[92][3]  ( .D(n1590), .CLK(clk_in), .RSTB(n7271), .Q(
        \FIFO[92][3] ) );
  DFFARX1 \FIFO_reg[92][2]  ( .D(n1589), .CLK(clk_in), .RSTB(n7271), .Q(
        \FIFO[92][2] ) );
  DFFARX1 \FIFO_reg[92][1]  ( .D(n1588), .CLK(clk_in), .RSTB(n7271), .Q(
        \FIFO[92][1] ) );
  DFFARX1 \FIFO_reg[92][0]  ( .D(n1587), .CLK(clk_in), .RSTB(n7271), .Q(
        \FIFO[92][0] ) );
  DFFARX1 \FIFO_reg[93][31]  ( .D(n1586), .CLK(clk_in), .RSTB(n7272), .Q(
        \FIFO[93][31] ) );
  DFFARX1 \FIFO_reg[93][30]  ( .D(n1585), .CLK(clk_in), .RSTB(n7272), .Q(
        \FIFO[93][30] ) );
  DFFARX1 \FIFO_reg[93][29]  ( .D(n1584), .CLK(clk_in), .RSTB(n7272), .Q(
        \FIFO[93][29] ) );
  DFFARX1 \FIFO_reg[93][28]  ( .D(n1583), .CLK(clk_in), .RSTB(n7272), .Q(
        \FIFO[93][28] ) );
  DFFARX1 \FIFO_reg[93][27]  ( .D(n1582), .CLK(clk_in), .RSTB(n7272), .Q(
        \FIFO[93][27] ) );
  DFFARX1 \FIFO_reg[93][26]  ( .D(n1581), .CLK(clk_in), .RSTB(n7272), .Q(
        \FIFO[93][26] ) );
  DFFARX1 \FIFO_reg[93][25]  ( .D(n1580), .CLK(clk_in), .RSTB(n7272), .Q(
        \FIFO[93][25] ) );
  DFFARX1 \FIFO_reg[93][24]  ( .D(n1579), .CLK(clk_in), .RSTB(n7272), .Q(
        \FIFO[93][24] ) );
  DFFARX1 \FIFO_reg[93][23]  ( .D(n1578), .CLK(clk_in), .RSTB(n7272), .Q(
        \FIFO[93][23] ) );
  DFFARX1 \FIFO_reg[93][22]  ( .D(n1577), .CLK(clk_in), .RSTB(n7272), .Q(
        \FIFO[93][22] ) );
  DFFARX1 \FIFO_reg[93][21]  ( .D(n1576), .CLK(clk_in), .RSTB(n7272), .Q(
        \FIFO[93][21] ) );
  DFFARX1 \FIFO_reg[93][20]  ( .D(n1575), .CLK(clk_in), .RSTB(n7272), .Q(
        \FIFO[93][20] ) );
  DFFARX1 \FIFO_reg[93][19]  ( .D(n1574), .CLK(clk_in), .RSTB(n7272), .Q(
        \FIFO[93][19] ) );
  DFFARX1 \FIFO_reg[93][18]  ( .D(n1573), .CLK(clk_in), .RSTB(n7272), .Q(
        \FIFO[93][18] ) );
  DFFARX1 \FIFO_reg[93][17]  ( .D(n1572), .CLK(clk_in), .RSTB(n7272), .Q(
        \FIFO[93][17] ) );
  DFFARX1 \FIFO_reg[93][16]  ( .D(n1571), .CLK(clk_in), .RSTB(n7272), .Q(
        \FIFO[93][16] ) );
  DFFARX1 \FIFO_reg[93][15]  ( .D(n1570), .CLK(clk_in), .RSTB(n7272), .Q(
        \FIFO[93][15] ) );
  DFFARX1 \FIFO_reg[93][14]  ( .D(n1569), .CLK(clk_in), .RSTB(n7272), .Q(
        \FIFO[93][14] ) );
  DFFARX1 \FIFO_reg[93][13]  ( .D(n1568), .CLK(clk_in), .RSTB(n7273), .Q(
        \FIFO[93][13] ) );
  DFFARX1 \FIFO_reg[93][12]  ( .D(n1567), .CLK(clk_in), .RSTB(n7273), .Q(
        \FIFO[93][12] ) );
  DFFARX1 \FIFO_reg[93][11]  ( .D(n1566), .CLK(clk_in), .RSTB(n7273), .Q(
        \FIFO[93][11] ) );
  DFFARX1 \FIFO_reg[93][10]  ( .D(n1565), .CLK(clk_in), .RSTB(n7273), .Q(
        \FIFO[93][10] ) );
  DFFARX1 \FIFO_reg[93][9]  ( .D(n1564), .CLK(clk_in), .RSTB(n7273), .Q(
        \FIFO[93][9] ) );
  DFFARX1 \FIFO_reg[93][8]  ( .D(n1563), .CLK(clk_in), .RSTB(n7273), .Q(
        \FIFO[93][8] ) );
  DFFARX1 \FIFO_reg[93][7]  ( .D(n1562), .CLK(clk_in), .RSTB(n7273), .Q(
        \FIFO[93][7] ) );
  DFFARX1 \FIFO_reg[93][6]  ( .D(n1561), .CLK(clk_in), .RSTB(n7273), .Q(
        \FIFO[93][6] ) );
  DFFARX1 \FIFO_reg[93][5]  ( .D(n1560), .CLK(clk_in), .RSTB(n7273), .Q(
        \FIFO[93][5] ) );
  DFFARX1 \FIFO_reg[93][4]  ( .D(n1559), .CLK(clk_in), .RSTB(n7273), .Q(
        \FIFO[93][4] ) );
  DFFARX1 \FIFO_reg[93][3]  ( .D(n1558), .CLK(clk_in), .RSTB(n7273), .Q(
        \FIFO[93][3] ) );
  DFFARX1 \FIFO_reg[93][2]  ( .D(n1557), .CLK(clk_in), .RSTB(n7273), .Q(
        \FIFO[93][2] ) );
  DFFARX1 \FIFO_reg[93][1]  ( .D(n1556), .CLK(clk_in), .RSTB(n7273), .Q(
        \FIFO[93][1] ) );
  DFFARX1 \FIFO_reg[93][0]  ( .D(n1555), .CLK(clk_in), .RSTB(n7273), .Q(
        \FIFO[93][0] ) );
  DFFARX1 \FIFO_reg[94][31]  ( .D(n1554), .CLK(clk_in), .RSTB(n7273), .Q(
        \FIFO[94][31] ) );
  DFFARX1 \FIFO_reg[94][30]  ( .D(n1553), .CLK(clk_in), .RSTB(n7273), .Q(
        \FIFO[94][30] ) );
  DFFARX1 \FIFO_reg[94][29]  ( .D(n1552), .CLK(clk_in), .RSTB(n7273), .Q(
        \FIFO[94][29] ) );
  DFFARX1 \FIFO_reg[94][28]  ( .D(n1551), .CLK(clk_in), .RSTB(n7273), .Q(
        \FIFO[94][28] ) );
  DFFARX1 \FIFO_reg[94][27]  ( .D(n1550), .CLK(clk_in), .RSTB(n7274), .Q(
        \FIFO[94][27] ) );
  DFFARX1 \FIFO_reg[94][26]  ( .D(n1549), .CLK(clk_in), .RSTB(n7274), .Q(
        \FIFO[94][26] ) );
  DFFARX1 \FIFO_reg[94][25]  ( .D(n1548), .CLK(clk_in), .RSTB(n7274), .Q(
        \FIFO[94][25] ) );
  DFFARX1 \FIFO_reg[94][24]  ( .D(n1547), .CLK(clk_in), .RSTB(n7274), .Q(
        \FIFO[94][24] ) );
  DFFARX1 \FIFO_reg[94][23]  ( .D(n1546), .CLK(clk_in), .RSTB(n7274), .Q(
        \FIFO[94][23] ) );
  DFFARX1 \FIFO_reg[94][22]  ( .D(n1545), .CLK(clk_in), .RSTB(n7274), .Q(
        \FIFO[94][22] ) );
  DFFARX1 \FIFO_reg[94][21]  ( .D(n1544), .CLK(clk_in), .RSTB(n7274), .Q(
        \FIFO[94][21] ) );
  DFFARX1 \FIFO_reg[94][20]  ( .D(n1543), .CLK(clk_in), .RSTB(n7274), .Q(
        \FIFO[94][20] ) );
  DFFARX1 \FIFO_reg[94][19]  ( .D(n1542), .CLK(clk_in), .RSTB(n7274), .Q(
        \FIFO[94][19] ) );
  DFFARX1 \FIFO_reg[94][18]  ( .D(n1541), .CLK(clk_in), .RSTB(n7274), .Q(
        \FIFO[94][18] ) );
  DFFARX1 \FIFO_reg[94][17]  ( .D(n1540), .CLK(clk_in), .RSTB(n7274), .Q(
        \FIFO[94][17] ) );
  DFFARX1 \FIFO_reg[94][16]  ( .D(n1539), .CLK(clk_in), .RSTB(n7274), .Q(
        \FIFO[94][16] ) );
  DFFARX1 \FIFO_reg[94][15]  ( .D(n1538), .CLK(clk_in), .RSTB(n7274), .Q(
        \FIFO[94][15] ) );
  DFFARX1 \FIFO_reg[94][14]  ( .D(n1537), .CLK(clk_in), .RSTB(n7274), .Q(
        \FIFO[94][14] ) );
  DFFARX1 \FIFO_reg[94][13]  ( .D(n1536), .CLK(clk_in), .RSTB(n7274), .Q(
        \FIFO[94][13] ) );
  DFFARX1 \FIFO_reg[94][12]  ( .D(n1535), .CLK(clk_in), .RSTB(n7274), .Q(
        \FIFO[94][12] ) );
  DFFARX1 \FIFO_reg[94][11]  ( .D(n1534), .CLK(clk_in), .RSTB(n7274), .Q(
        \FIFO[94][11] ) );
  DFFARX1 \FIFO_reg[94][10]  ( .D(n1533), .CLK(clk_in), .RSTB(n7274), .Q(
        \FIFO[94][10] ) );
  DFFARX1 \FIFO_reg[94][9]  ( .D(n1532), .CLK(clk_in), .RSTB(n7275), .Q(
        \FIFO[94][9] ) );
  DFFARX1 \FIFO_reg[94][8]  ( .D(n1531), .CLK(clk_in), .RSTB(n7275), .Q(
        \FIFO[94][8] ) );
  DFFARX1 \FIFO_reg[94][7]  ( .D(n1530), .CLK(clk_in), .RSTB(n7275), .Q(
        \FIFO[94][7] ) );
  DFFARX1 \FIFO_reg[94][6]  ( .D(n1529), .CLK(clk_in), .RSTB(n7275), .Q(
        \FIFO[94][6] ) );
  DFFARX1 \FIFO_reg[94][5]  ( .D(n1528), .CLK(clk_in), .RSTB(n7275), .Q(
        \FIFO[94][5] ) );
  DFFARX1 \FIFO_reg[94][4]  ( .D(n1527), .CLK(clk_in), .RSTB(n7275), .Q(
        \FIFO[94][4] ) );
  DFFARX1 \FIFO_reg[94][3]  ( .D(n1526), .CLK(clk_in), .RSTB(n7275), .Q(
        \FIFO[94][3] ) );
  DFFARX1 \FIFO_reg[94][2]  ( .D(n1525), .CLK(clk_in), .RSTB(n7275), .Q(
        \FIFO[94][2] ) );
  DFFARX1 \FIFO_reg[94][1]  ( .D(n1524), .CLK(clk_in), .RSTB(n7275), .Q(
        \FIFO[94][1] ) );
  DFFARX1 \FIFO_reg[94][0]  ( .D(n1523), .CLK(clk_in), .RSTB(n7275), .Q(
        \FIFO[94][0] ) );
  DFFARX1 \FIFO_reg[95][31]  ( .D(n1522), .CLK(clk_in), .RSTB(n7275), .Q(
        \FIFO[95][31] ) );
  DFFARX1 \FIFO_reg[95][30]  ( .D(n1521), .CLK(clk_in), .RSTB(n7275), .Q(
        \FIFO[95][30] ) );
  DFFARX1 \FIFO_reg[95][29]  ( .D(n1520), .CLK(clk_in), .RSTB(n7275), .Q(
        \FIFO[95][29] ) );
  DFFARX1 \FIFO_reg[95][28]  ( .D(n1519), .CLK(clk_in), .RSTB(n7275), .Q(
        \FIFO[95][28] ) );
  DFFARX1 \FIFO_reg[95][27]  ( .D(n1518), .CLK(clk_in), .RSTB(n7275), .Q(
        \FIFO[95][27] ) );
  DFFARX1 \FIFO_reg[95][26]  ( .D(n1517), .CLK(clk_in), .RSTB(n7275), .Q(
        \FIFO[95][26] ) );
  DFFARX1 \FIFO_reg[95][25]  ( .D(n1516), .CLK(clk_in), .RSTB(n7275), .Q(
        \FIFO[95][25] ) );
  DFFARX1 \FIFO_reg[95][24]  ( .D(n1515), .CLK(clk_in), .RSTB(n7275), .Q(
        \FIFO[95][24] ) );
  DFFARX1 \FIFO_reg[95][23]  ( .D(n1514), .CLK(clk_in), .RSTB(n7276), .Q(
        \FIFO[95][23] ) );
  DFFARX1 \FIFO_reg[95][22]  ( .D(n1513), .CLK(clk_in), .RSTB(n7276), .Q(
        \FIFO[95][22] ) );
  DFFARX1 \FIFO_reg[95][21]  ( .D(n1512), .CLK(clk_in), .RSTB(n7276), .Q(
        \FIFO[95][21] ) );
  DFFARX1 \FIFO_reg[95][20]  ( .D(n1511), .CLK(clk_in), .RSTB(n7276), .Q(
        \FIFO[95][20] ) );
  DFFARX1 \FIFO_reg[95][19]  ( .D(n1510), .CLK(clk_in), .RSTB(n7276), .Q(
        \FIFO[95][19] ) );
  DFFARX1 \FIFO_reg[95][18]  ( .D(n1509), .CLK(clk_in), .RSTB(n7276), .Q(
        \FIFO[95][18] ) );
  DFFARX1 \FIFO_reg[95][17]  ( .D(n1508), .CLK(clk_in), .RSTB(n7276), .Q(
        \FIFO[95][17] ) );
  DFFARX1 \FIFO_reg[95][16]  ( .D(n1507), .CLK(clk_in), .RSTB(n7276), .Q(
        \FIFO[95][16] ) );
  DFFARX1 \FIFO_reg[95][15]  ( .D(n1506), .CLK(clk_in), .RSTB(n7276), .Q(
        \FIFO[95][15] ) );
  DFFARX1 \FIFO_reg[95][14]  ( .D(n1505), .CLK(clk_in), .RSTB(n7276), .Q(
        \FIFO[95][14] ) );
  DFFARX1 \FIFO_reg[95][13]  ( .D(n1504), .CLK(clk_in), .RSTB(n7276), .Q(
        \FIFO[95][13] ) );
  DFFARX1 \FIFO_reg[95][12]  ( .D(n1503), .CLK(clk_in), .RSTB(n7276), .Q(
        \FIFO[95][12] ) );
  DFFARX1 \FIFO_reg[95][11]  ( .D(n1502), .CLK(clk_in), .RSTB(n7276), .Q(
        \FIFO[95][11] ) );
  DFFARX1 \FIFO_reg[95][10]  ( .D(n1501), .CLK(clk_in), .RSTB(n7276), .Q(
        \FIFO[95][10] ) );
  DFFARX1 \FIFO_reg[95][9]  ( .D(n1500), .CLK(clk_in), .RSTB(n7276), .Q(
        \FIFO[95][9] ) );
  DFFARX1 \FIFO_reg[95][8]  ( .D(n1499), .CLK(clk_in), .RSTB(n7276), .Q(
        \FIFO[95][8] ) );
  DFFARX1 \FIFO_reg[95][7]  ( .D(n1498), .CLK(clk_in), .RSTB(n7276), .Q(
        \FIFO[95][7] ) );
  DFFARX1 \FIFO_reg[95][6]  ( .D(n1497), .CLK(clk_in), .RSTB(n7276), .Q(
        \FIFO[95][6] ) );
  DFFARX1 \FIFO_reg[95][5]  ( .D(n1496), .CLK(clk_in), .RSTB(n7277), .Q(
        \FIFO[95][5] ) );
  DFFARX1 \FIFO_reg[95][4]  ( .D(n1495), .CLK(clk_in), .RSTB(n7277), .Q(
        \FIFO[95][4] ) );
  DFFARX1 \FIFO_reg[95][3]  ( .D(n1494), .CLK(clk_in), .RSTB(n7277), .Q(
        \FIFO[95][3] ) );
  DFFARX1 \FIFO_reg[95][2]  ( .D(n1493), .CLK(clk_in), .RSTB(n7277), .Q(
        \FIFO[95][2] ) );
  DFFARX1 \FIFO_reg[95][1]  ( .D(n1492), .CLK(clk_in), .RSTB(n7277), .Q(
        \FIFO[95][1] ) );
  DFFARX1 \FIFO_reg[95][0]  ( .D(n1491), .CLK(clk_in), .RSTB(n7277), .Q(
        \FIFO[95][0] ) );
  DFFARX1 \FIFO_reg[96][31]  ( .D(n1490), .CLK(clk_in), .RSTB(n7277), .Q(
        \FIFO[96][31] ) );
  DFFARX1 \FIFO_reg[96][30]  ( .D(n1489), .CLK(clk_in), .RSTB(n7277), .Q(
        \FIFO[96][30] ) );
  DFFARX1 \FIFO_reg[96][29]  ( .D(n1488), .CLK(clk_in), .RSTB(n7277), .Q(
        \FIFO[96][29] ) );
  DFFARX1 \FIFO_reg[96][28]  ( .D(n1487), .CLK(clk_in), .RSTB(n7277), .Q(
        \FIFO[96][28] ) );
  DFFARX1 \FIFO_reg[96][27]  ( .D(n1486), .CLK(clk_in), .RSTB(n7277), .Q(
        \FIFO[96][27] ) );
  DFFARX1 \FIFO_reg[96][26]  ( .D(n1485), .CLK(clk_in), .RSTB(n7277), .Q(
        \FIFO[96][26] ) );
  DFFARX1 \FIFO_reg[96][25]  ( .D(n1484), .CLK(clk_in), .RSTB(n7277), .Q(
        \FIFO[96][25] ) );
  DFFARX1 \FIFO_reg[96][24]  ( .D(n1483), .CLK(clk_in), .RSTB(n7277), .Q(
        \FIFO[96][24] ) );
  DFFARX1 \FIFO_reg[96][23]  ( .D(n1482), .CLK(clk_in), .RSTB(n7277), .Q(
        \FIFO[96][23] ) );
  DFFARX1 \FIFO_reg[96][22]  ( .D(n1481), .CLK(clk_in), .RSTB(n7277), .Q(
        \FIFO[96][22] ) );
  DFFARX1 \FIFO_reg[96][21]  ( .D(n1480), .CLK(clk_in), .RSTB(n7277), .Q(
        \FIFO[96][21] ) );
  DFFARX1 \FIFO_reg[96][20]  ( .D(n1479), .CLK(clk_in), .RSTB(n7277), .Q(
        \FIFO[96][20] ) );
  DFFARX1 \FIFO_reg[96][19]  ( .D(n1478), .CLK(clk_in), .RSTB(n7278), .Q(
        \FIFO[96][19] ) );
  DFFARX1 \FIFO_reg[96][18]  ( .D(n1477), .CLK(clk_in), .RSTB(n7278), .Q(
        \FIFO[96][18] ) );
  DFFARX1 \FIFO_reg[96][17]  ( .D(n1476), .CLK(clk_in), .RSTB(n7278), .Q(
        \FIFO[96][17] ) );
  DFFARX1 \FIFO_reg[96][16]  ( .D(n1475), .CLK(clk_in), .RSTB(n7278), .Q(
        \FIFO[96][16] ) );
  DFFARX1 \FIFO_reg[96][15]  ( .D(n1474), .CLK(clk_in), .RSTB(n7278), .Q(
        \FIFO[96][15] ) );
  DFFARX1 \FIFO_reg[96][14]  ( .D(n1473), .CLK(clk_in), .RSTB(n7278), .Q(
        \FIFO[96][14] ) );
  DFFARX1 \FIFO_reg[96][13]  ( .D(n1472), .CLK(clk_in), .RSTB(n7278), .Q(
        \FIFO[96][13] ) );
  DFFARX1 \FIFO_reg[96][12]  ( .D(n1471), .CLK(clk_in), .RSTB(n7278), .Q(
        \FIFO[96][12] ) );
  DFFARX1 \FIFO_reg[96][11]  ( .D(n1470), .CLK(clk_in), .RSTB(n7278), .Q(
        \FIFO[96][11] ) );
  DFFARX1 \FIFO_reg[96][10]  ( .D(n1469), .CLK(clk_in), .RSTB(n7278), .Q(
        \FIFO[96][10] ) );
  DFFARX1 \FIFO_reg[96][9]  ( .D(n1468), .CLK(clk_in), .RSTB(n7278), .Q(
        \FIFO[96][9] ) );
  DFFARX1 \FIFO_reg[96][8]  ( .D(n1467), .CLK(clk_in), .RSTB(n7278), .Q(
        \FIFO[96][8] ) );
  DFFARX1 \FIFO_reg[96][7]  ( .D(n1466), .CLK(clk_in), .RSTB(n7278), .Q(
        \FIFO[96][7] ) );
  DFFARX1 \FIFO_reg[96][6]  ( .D(n1465), .CLK(clk_in), .RSTB(n7278), .Q(
        \FIFO[96][6] ) );
  DFFARX1 \FIFO_reg[96][5]  ( .D(n1464), .CLK(clk_in), .RSTB(n7278), .Q(
        \FIFO[96][5] ) );
  DFFARX1 \FIFO_reg[96][4]  ( .D(n1463), .CLK(clk_in), .RSTB(n7278), .Q(
        \FIFO[96][4] ) );
  DFFARX1 \FIFO_reg[96][3]  ( .D(n1462), .CLK(clk_in), .RSTB(n7278), .Q(
        \FIFO[96][3] ) );
  DFFARX1 \FIFO_reg[96][2]  ( .D(n1461), .CLK(clk_in), .RSTB(n7278), .Q(
        \FIFO[96][2] ) );
  DFFARX1 \FIFO_reg[96][1]  ( .D(n1460), .CLK(clk_in), .RSTB(n7279), .Q(
        \FIFO[96][1] ) );
  DFFARX1 \FIFO_reg[96][0]  ( .D(n1459), .CLK(clk_in), .RSTB(n7279), .Q(
        \FIFO[96][0] ) );
  DFFARX1 \FIFO_reg[97][31]  ( .D(n1458), .CLK(clk_in), .RSTB(n7279), .Q(
        \FIFO[97][31] ) );
  DFFARX1 \FIFO_reg[97][30]  ( .D(n1457), .CLK(clk_in), .RSTB(n7279), .Q(
        \FIFO[97][30] ) );
  DFFARX1 \FIFO_reg[97][29]  ( .D(n1456), .CLK(clk_in), .RSTB(n7279), .Q(
        \FIFO[97][29] ) );
  DFFARX1 \FIFO_reg[97][28]  ( .D(n1455), .CLK(clk_in), .RSTB(n7279), .Q(
        \FIFO[97][28] ) );
  DFFARX1 \FIFO_reg[97][27]  ( .D(n1454), .CLK(clk_in), .RSTB(n7279), .Q(
        \FIFO[97][27] ) );
  DFFARX1 \FIFO_reg[97][26]  ( .D(n1453), .CLK(clk_in), .RSTB(n7279), .Q(
        \FIFO[97][26] ) );
  DFFARX1 \FIFO_reg[97][25]  ( .D(n1452), .CLK(clk_in), .RSTB(n7279), .Q(
        \FIFO[97][25] ) );
  DFFARX1 \FIFO_reg[97][24]  ( .D(n1451), .CLK(clk_in), .RSTB(n7279), .Q(
        \FIFO[97][24] ) );
  DFFARX1 \FIFO_reg[97][23]  ( .D(n1450), .CLK(clk_in), .RSTB(n7279), .Q(
        \FIFO[97][23] ) );
  DFFARX1 \FIFO_reg[97][22]  ( .D(n1449), .CLK(clk_in), .RSTB(n7279), .Q(
        \FIFO[97][22] ) );
  DFFARX1 \FIFO_reg[97][21]  ( .D(n1448), .CLK(clk_in), .RSTB(n7279), .Q(
        \FIFO[97][21] ) );
  DFFARX1 \FIFO_reg[97][20]  ( .D(n1447), .CLK(clk_in), .RSTB(n7279), .Q(
        \FIFO[97][20] ) );
  DFFARX1 \FIFO_reg[97][19]  ( .D(n1446), .CLK(clk_in), .RSTB(n7279), .Q(
        \FIFO[97][19] ) );
  DFFARX1 \FIFO_reg[97][18]  ( .D(n1445), .CLK(clk_in), .RSTB(n7279), .Q(
        \FIFO[97][18] ) );
  DFFARX1 \FIFO_reg[97][17]  ( .D(n1444), .CLK(clk_in), .RSTB(n7279), .Q(
        \FIFO[97][17] ) );
  DFFARX1 \FIFO_reg[97][16]  ( .D(n1443), .CLK(clk_in), .RSTB(n7279), .Q(
        \FIFO[97][16] ) );
  DFFARX1 \FIFO_reg[97][15]  ( .D(n1442), .CLK(clk_in), .RSTB(n7280), .Q(
        \FIFO[97][15] ) );
  DFFARX1 \FIFO_reg[97][14]  ( .D(n1441), .CLK(clk_in), .RSTB(n7280), .Q(
        \FIFO[97][14] ) );
  DFFARX1 \FIFO_reg[97][13]  ( .D(n1440), .CLK(clk_in), .RSTB(n7280), .Q(
        \FIFO[97][13] ) );
  DFFARX1 \FIFO_reg[97][12]  ( .D(n1439), .CLK(clk_in), .RSTB(n7280), .Q(
        \FIFO[97][12] ) );
  DFFARX1 \FIFO_reg[97][11]  ( .D(n1438), .CLK(clk_in), .RSTB(n7280), .Q(
        \FIFO[97][11] ) );
  DFFARX1 \FIFO_reg[97][10]  ( .D(n1437), .CLK(clk_in), .RSTB(n7280), .Q(
        \FIFO[97][10] ) );
  DFFARX1 \FIFO_reg[97][9]  ( .D(n1436), .CLK(clk_in), .RSTB(n7280), .Q(
        \FIFO[97][9] ) );
  DFFARX1 \FIFO_reg[97][8]  ( .D(n1435), .CLK(clk_in), .RSTB(n7280), .Q(
        \FIFO[97][8] ) );
  DFFARX1 \FIFO_reg[97][7]  ( .D(n1434), .CLK(clk_in), .RSTB(n7280), .Q(
        \FIFO[97][7] ) );
  DFFARX1 \FIFO_reg[97][6]  ( .D(n1433), .CLK(clk_in), .RSTB(n7280), .Q(
        \FIFO[97][6] ) );
  DFFARX1 \FIFO_reg[97][5]  ( .D(n1432), .CLK(clk_in), .RSTB(n7280), .Q(
        \FIFO[97][5] ) );
  DFFARX1 \FIFO_reg[97][4]  ( .D(n1431), .CLK(clk_in), .RSTB(n7280), .Q(
        \FIFO[97][4] ) );
  DFFARX1 \FIFO_reg[97][3]  ( .D(n1430), .CLK(clk_in), .RSTB(n7280), .Q(
        \FIFO[97][3] ) );
  DFFARX1 \FIFO_reg[97][2]  ( .D(n1429), .CLK(clk_in), .RSTB(n7280), .Q(
        \FIFO[97][2] ) );
  DFFARX1 \FIFO_reg[97][1]  ( .D(n1428), .CLK(clk_in), .RSTB(n7280), .Q(
        \FIFO[97][1] ) );
  DFFARX1 \FIFO_reg[97][0]  ( .D(n1427), .CLK(clk_in), .RSTB(n7280), .Q(
        \FIFO[97][0] ) );
  DFFARX1 \FIFO_reg[98][31]  ( .D(n1426), .CLK(clk_in), .RSTB(n7280), .Q(
        \FIFO[98][31] ) );
  DFFARX1 \FIFO_reg[98][30]  ( .D(n1425), .CLK(clk_in), .RSTB(n7280), .Q(
        \FIFO[98][30] ) );
  DFFARX1 \FIFO_reg[98][29]  ( .D(n1424), .CLK(clk_in), .RSTB(n7281), .Q(
        \FIFO[98][29] ) );
  DFFARX1 \FIFO_reg[98][28]  ( .D(n1423), .CLK(clk_in), .RSTB(n7281), .Q(
        \FIFO[98][28] ) );
  DFFARX1 \FIFO_reg[98][27]  ( .D(n1422), .CLK(clk_in), .RSTB(n7281), .Q(
        \FIFO[98][27] ) );
  DFFARX1 \FIFO_reg[98][26]  ( .D(n1421), .CLK(clk_in), .RSTB(n7281), .Q(
        \FIFO[98][26] ) );
  DFFARX1 \FIFO_reg[98][25]  ( .D(n1420), .CLK(clk_in), .RSTB(n7281), .Q(
        \FIFO[98][25] ) );
  DFFARX1 \FIFO_reg[98][24]  ( .D(n1419), .CLK(clk_in), .RSTB(n7281), .Q(
        \FIFO[98][24] ) );
  DFFARX1 \FIFO_reg[98][23]  ( .D(n1418), .CLK(clk_in), .RSTB(n7281), .Q(
        \FIFO[98][23] ) );
  DFFARX1 \FIFO_reg[98][22]  ( .D(n1417), .CLK(clk_in), .RSTB(n7281), .Q(
        \FIFO[98][22] ) );
  DFFARX1 \FIFO_reg[98][21]  ( .D(n1416), .CLK(clk_in), .RSTB(n7281), .Q(
        \FIFO[98][21] ) );
  DFFARX1 \FIFO_reg[98][20]  ( .D(n1415), .CLK(clk_in), .RSTB(n7281), .Q(
        \FIFO[98][20] ) );
  DFFARX1 \FIFO_reg[98][19]  ( .D(n1414), .CLK(clk_in), .RSTB(n7281), .Q(
        \FIFO[98][19] ) );
  DFFARX1 \FIFO_reg[98][18]  ( .D(n1413), .CLK(clk_in), .RSTB(n7281), .Q(
        \FIFO[98][18] ) );
  DFFARX1 \FIFO_reg[98][17]  ( .D(n1412), .CLK(clk_in), .RSTB(n7281), .Q(
        \FIFO[98][17] ) );
  DFFARX1 \FIFO_reg[98][16]  ( .D(n1411), .CLK(clk_in), .RSTB(n7281), .Q(
        \FIFO[98][16] ) );
  DFFARX1 \FIFO_reg[98][15]  ( .D(n1410), .CLK(clk_in), .RSTB(n7281), .Q(
        \FIFO[98][15] ) );
  DFFARX1 \FIFO_reg[98][14]  ( .D(n1409), .CLK(clk_in), .RSTB(n7281), .Q(
        \FIFO[98][14] ) );
  DFFARX1 \FIFO_reg[98][13]  ( .D(n1408), .CLK(clk_in), .RSTB(n7281), .Q(
        \FIFO[98][13] ) );
  DFFARX1 \FIFO_reg[98][12]  ( .D(n1407), .CLK(clk_in), .RSTB(n7281), .Q(
        \FIFO[98][12] ) );
  DFFARX1 \FIFO_reg[98][11]  ( .D(n1406), .CLK(clk_in), .RSTB(n7282), .Q(
        \FIFO[98][11] ) );
  DFFARX1 \FIFO_reg[98][10]  ( .D(n1405), .CLK(clk_in), .RSTB(n7282), .Q(
        \FIFO[98][10] ) );
  DFFARX1 \FIFO_reg[98][9]  ( .D(n1404), .CLK(clk_in), .RSTB(n7282), .Q(
        \FIFO[98][9] ) );
  DFFARX1 \FIFO_reg[98][8]  ( .D(n1403), .CLK(clk_in), .RSTB(n7282), .Q(
        \FIFO[98][8] ) );
  DFFARX1 \FIFO_reg[98][7]  ( .D(n1402), .CLK(clk_in), .RSTB(n7282), .Q(
        \FIFO[98][7] ) );
  DFFARX1 \FIFO_reg[98][6]  ( .D(n1401), .CLK(clk_in), .RSTB(n7282), .Q(
        \FIFO[98][6] ) );
  DFFARX1 \FIFO_reg[98][5]  ( .D(n1400), .CLK(clk_in), .RSTB(n7282), .Q(
        \FIFO[98][5] ) );
  DFFARX1 \FIFO_reg[98][4]  ( .D(n1399), .CLK(clk_in), .RSTB(n7282), .Q(
        \FIFO[98][4] ) );
  DFFARX1 \FIFO_reg[98][3]  ( .D(n1398), .CLK(clk_in), .RSTB(n7282), .Q(
        \FIFO[98][3] ) );
  DFFARX1 \FIFO_reg[98][2]  ( .D(n1397), .CLK(clk_in), .RSTB(n7282), .Q(
        \FIFO[98][2] ) );
  DFFARX1 \FIFO_reg[98][1]  ( .D(n1396), .CLK(clk_in), .RSTB(n7282), .Q(
        \FIFO[98][1] ) );
  DFFARX1 \FIFO_reg[98][0]  ( .D(n1395), .CLK(clk_in), .RSTB(n7282), .Q(
        \FIFO[98][0] ) );
  DFFARX1 \FIFO_reg[99][31]  ( .D(n1394), .CLK(clk_in), .RSTB(n7282), .Q(
        \FIFO[99][31] ) );
  DFFARX1 \FIFO_reg[99][30]  ( .D(n1393), .CLK(clk_in), .RSTB(n7282), .Q(
        \FIFO[99][30] ) );
  DFFARX1 \FIFO_reg[99][29]  ( .D(n1392), .CLK(clk_in), .RSTB(n7282), .Q(
        \FIFO[99][29] ) );
  DFFARX1 \FIFO_reg[99][28]  ( .D(n1391), .CLK(clk_in), .RSTB(n7282), .Q(
        \FIFO[99][28] ) );
  DFFARX1 \FIFO_reg[99][27]  ( .D(n1390), .CLK(clk_in), .RSTB(n7282), .Q(
        \FIFO[99][27] ) );
  DFFARX1 \FIFO_reg[99][26]  ( .D(n1389), .CLK(clk_in), .RSTB(n7282), .Q(
        \FIFO[99][26] ) );
  DFFARX1 \FIFO_reg[99][25]  ( .D(n1388), .CLK(clk_in), .RSTB(n7283), .Q(
        \FIFO[99][25] ) );
  DFFARX1 \FIFO_reg[99][24]  ( .D(n1387), .CLK(clk_in), .RSTB(n7283), .Q(
        \FIFO[99][24] ) );
  DFFARX1 \FIFO_reg[99][23]  ( .D(n1386), .CLK(clk_in), .RSTB(n7283), .Q(
        \FIFO[99][23] ) );
  DFFARX1 \FIFO_reg[99][22]  ( .D(n1385), .CLK(clk_in), .RSTB(n7283), .Q(
        \FIFO[99][22] ) );
  DFFARX1 \FIFO_reg[99][21]  ( .D(n1384), .CLK(clk_in), .RSTB(n7283), .Q(
        \FIFO[99][21] ) );
  DFFARX1 \FIFO_reg[99][20]  ( .D(n1383), .CLK(clk_in), .RSTB(n7283), .Q(
        \FIFO[99][20] ) );
  DFFARX1 \FIFO_reg[99][19]  ( .D(n1382), .CLK(clk_in), .RSTB(n7283), .Q(
        \FIFO[99][19] ) );
  DFFARX1 \FIFO_reg[99][18]  ( .D(n1381), .CLK(clk_in), .RSTB(n7283), .Q(
        \FIFO[99][18] ) );
  DFFARX1 \FIFO_reg[99][17]  ( .D(n1380), .CLK(clk_in), .RSTB(n7283), .Q(
        \FIFO[99][17] ) );
  DFFARX1 \FIFO_reg[99][16]  ( .D(n1379), .CLK(clk_in), .RSTB(n7283), .Q(
        \FIFO[99][16] ) );
  DFFARX1 \FIFO_reg[99][15]  ( .D(n1378), .CLK(clk_in), .RSTB(n7283), .Q(
        \FIFO[99][15] ) );
  DFFARX1 \FIFO_reg[99][14]  ( .D(n1377), .CLK(clk_in), .RSTB(n7283), .Q(
        \FIFO[99][14] ) );
  DFFARX1 \FIFO_reg[99][13]  ( .D(n1376), .CLK(clk_in), .RSTB(n7283), .Q(
        \FIFO[99][13] ) );
  DFFARX1 \FIFO_reg[99][12]  ( .D(n1375), .CLK(clk_in), .RSTB(n7283), .Q(
        \FIFO[99][12] ) );
  DFFARX1 \FIFO_reg[99][11]  ( .D(n1374), .CLK(clk_in), .RSTB(n7283), .Q(
        \FIFO[99][11] ) );
  DFFARX1 \FIFO_reg[99][10]  ( .D(n1373), .CLK(clk_in), .RSTB(n7283), .Q(
        \FIFO[99][10] ) );
  DFFARX1 \FIFO_reg[99][9]  ( .D(n1372), .CLK(clk_in), .RSTB(n7283), .Q(
        \FIFO[99][9] ) );
  DFFARX1 \FIFO_reg[99][8]  ( .D(n1371), .CLK(clk_in), .RSTB(n7283), .Q(
        \FIFO[99][8] ) );
  DFFARX1 \FIFO_reg[99][7]  ( .D(n1370), .CLK(clk_in), .RSTB(n7284), .Q(
        \FIFO[99][7] ) );
  DFFARX1 \FIFO_reg[99][6]  ( .D(n1369), .CLK(clk_in), .RSTB(n7284), .Q(
        \FIFO[99][6] ) );
  DFFARX1 \FIFO_reg[99][5]  ( .D(n1368), .CLK(clk_in), .RSTB(n7284), .Q(
        \FIFO[99][5] ) );
  DFFARX1 \FIFO_reg[99][4]  ( .D(n1367), .CLK(clk_in), .RSTB(n7284), .Q(
        \FIFO[99][4] ) );
  DFFARX1 \FIFO_reg[99][3]  ( .D(n1366), .CLK(clk_in), .RSTB(n7284), .Q(
        \FIFO[99][3] ) );
  DFFARX1 \FIFO_reg[99][2]  ( .D(n1365), .CLK(clk_in), .RSTB(n7284), .Q(
        \FIFO[99][2] ) );
  DFFARX1 \FIFO_reg[99][1]  ( .D(n1364), .CLK(clk_in), .RSTB(n7284), .Q(
        \FIFO[99][1] ) );
  DFFARX1 \FIFO_reg[99][0]  ( .D(n1363), .CLK(clk_in), .RSTB(n7284), .Q(
        \FIFO[99][0] ) );
  DFFARX1 \FIFO_reg[100][31]  ( .D(n1362), .CLK(clk_in), .RSTB(n7284), .Q(
        \FIFO[100][31] ) );
  DFFARX1 \FIFO_reg[100][30]  ( .D(n1361), .CLK(clk_in), .RSTB(n7284), .Q(
        \FIFO[100][30] ) );
  DFFARX1 \FIFO_reg[100][29]  ( .D(n1360), .CLK(clk_in), .RSTB(n7284), .Q(
        \FIFO[100][29] ) );
  DFFARX1 \FIFO_reg[100][28]  ( .D(n1359), .CLK(clk_in), .RSTB(n7284), .Q(
        \FIFO[100][28] ) );
  DFFARX1 \FIFO_reg[100][27]  ( .D(n1358), .CLK(clk_in), .RSTB(n7284), .Q(
        \FIFO[100][27] ) );
  DFFARX1 \FIFO_reg[100][26]  ( .D(n1357), .CLK(clk_in), .RSTB(n7284), .Q(
        \FIFO[100][26] ) );
  DFFARX1 \FIFO_reg[100][25]  ( .D(n1356), .CLK(clk_in), .RSTB(n7284), .Q(
        \FIFO[100][25] ) );
  DFFARX1 \FIFO_reg[100][24]  ( .D(n1355), .CLK(clk_in), .RSTB(n7284), .Q(
        \FIFO[100][24] ) );
  DFFARX1 \FIFO_reg[100][23]  ( .D(n1354), .CLK(clk_in), .RSTB(n7284), .Q(
        \FIFO[100][23] ) );
  DFFARX1 \FIFO_reg[100][22]  ( .D(n1353), .CLK(clk_in), .RSTB(n7284), .Q(
        \FIFO[100][22] ) );
  DFFARX1 \FIFO_reg[100][21]  ( .D(n1352), .CLK(clk_in), .RSTB(n7285), .Q(
        \FIFO[100][21] ) );
  DFFARX1 \FIFO_reg[100][20]  ( .D(n1351), .CLK(clk_in), .RSTB(n7285), .Q(
        \FIFO[100][20] ) );
  DFFARX1 \FIFO_reg[100][19]  ( .D(n1350), .CLK(clk_in), .RSTB(n7285), .Q(
        \FIFO[100][19] ) );
  DFFARX1 \FIFO_reg[100][18]  ( .D(n1349), .CLK(clk_in), .RSTB(n7285), .Q(
        \FIFO[100][18] ) );
  DFFARX1 \FIFO_reg[100][17]  ( .D(n1348), .CLK(clk_in), .RSTB(n7285), .Q(
        \FIFO[100][17] ) );
  DFFARX1 \FIFO_reg[100][16]  ( .D(n1347), .CLK(clk_in), .RSTB(n7285), .Q(
        \FIFO[100][16] ) );
  DFFARX1 \FIFO_reg[100][15]  ( .D(n1346), .CLK(clk_in), .RSTB(n7285), .Q(
        \FIFO[100][15] ) );
  DFFARX1 \FIFO_reg[100][14]  ( .D(n1345), .CLK(clk_in), .RSTB(n7285), .Q(
        \FIFO[100][14] ) );
  DFFARX1 \FIFO_reg[100][13]  ( .D(n1344), .CLK(clk_in), .RSTB(n7285), .Q(
        \FIFO[100][13] ) );
  DFFARX1 \FIFO_reg[100][12]  ( .D(n1343), .CLK(clk_in), .RSTB(n7285), .Q(
        \FIFO[100][12] ) );
  DFFARX1 \FIFO_reg[100][11]  ( .D(n1342), .CLK(clk_in), .RSTB(n7285), .Q(
        \FIFO[100][11] ) );
  DFFARX1 \FIFO_reg[100][10]  ( .D(n1341), .CLK(clk_in), .RSTB(n7285), .Q(
        \FIFO[100][10] ) );
  DFFARX1 \FIFO_reg[100][9]  ( .D(n1340), .CLK(clk_in), .RSTB(n7285), .Q(
        \FIFO[100][9] ) );
  DFFARX1 \FIFO_reg[100][8]  ( .D(n1339), .CLK(clk_in), .RSTB(n7285), .Q(
        \FIFO[100][8] ) );
  DFFARX1 \FIFO_reg[100][7]  ( .D(n1338), .CLK(clk_in), .RSTB(n7285), .Q(
        \FIFO[100][7] ) );
  DFFARX1 \FIFO_reg[100][6]  ( .D(n1337), .CLK(clk_in), .RSTB(n7285), .Q(
        \FIFO[100][6] ) );
  DFFARX1 \FIFO_reg[100][5]  ( .D(n1336), .CLK(clk_in), .RSTB(n7285), .Q(
        \FIFO[100][5] ) );
  DFFARX1 \FIFO_reg[100][4]  ( .D(n1335), .CLK(clk_in), .RSTB(n7285), .Q(
        \FIFO[100][4] ) );
  DFFARX1 \FIFO_reg[100][3]  ( .D(n1334), .CLK(clk_in), .RSTB(n7286), .Q(
        \FIFO[100][3] ) );
  DFFARX1 \FIFO_reg[100][2]  ( .D(n1333), .CLK(clk_in), .RSTB(n7286), .Q(
        \FIFO[100][2] ) );
  DFFARX1 \FIFO_reg[100][1]  ( .D(n1332), .CLK(clk_in), .RSTB(n7286), .Q(
        \FIFO[100][1] ) );
  DFFARX1 \FIFO_reg[100][0]  ( .D(n1331), .CLK(clk_in), .RSTB(n7286), .Q(
        \FIFO[100][0] ) );
  DFFARX1 \FIFO_reg[101][31]  ( .D(n1330), .CLK(clk_in), .RSTB(n7286), .Q(
        \FIFO[101][31] ) );
  DFFARX1 \FIFO_reg[101][30]  ( .D(n1329), .CLK(clk_in), .RSTB(n7286), .Q(
        \FIFO[101][30] ) );
  DFFARX1 \FIFO_reg[101][29]  ( .D(n1328), .CLK(clk_in), .RSTB(n7286), .Q(
        \FIFO[101][29] ) );
  DFFARX1 \FIFO_reg[101][28]  ( .D(n1327), .CLK(clk_in), .RSTB(n7286), .Q(
        \FIFO[101][28] ) );
  DFFARX1 \FIFO_reg[101][27]  ( .D(n1326), .CLK(clk_in), .RSTB(n7286), .Q(
        \FIFO[101][27] ) );
  DFFARX1 \FIFO_reg[101][26]  ( .D(n1325), .CLK(clk_in), .RSTB(n7286), .Q(
        \FIFO[101][26] ) );
  DFFARX1 \FIFO_reg[101][25]  ( .D(n1324), .CLK(clk_in), .RSTB(n7286), .Q(
        \FIFO[101][25] ) );
  DFFARX1 \FIFO_reg[101][24]  ( .D(n1323), .CLK(clk_in), .RSTB(n7286), .Q(
        \FIFO[101][24] ) );
  DFFARX1 \FIFO_reg[101][23]  ( .D(n1322), .CLK(clk_in), .RSTB(n7286), .Q(
        \FIFO[101][23] ) );
  DFFARX1 \FIFO_reg[101][22]  ( .D(n1321), .CLK(clk_in), .RSTB(n7286), .Q(
        \FIFO[101][22] ) );
  DFFARX1 \FIFO_reg[101][21]  ( .D(n1320), .CLK(clk_in), .RSTB(n7286), .Q(
        \FIFO[101][21] ) );
  DFFARX1 \FIFO_reg[101][20]  ( .D(n1319), .CLK(clk_in), .RSTB(n7286), .Q(
        \FIFO[101][20] ) );
  DFFARX1 \FIFO_reg[101][19]  ( .D(n1318), .CLK(clk_in), .RSTB(n7286), .Q(
        \FIFO[101][19] ) );
  DFFARX1 \FIFO_reg[101][18]  ( .D(n1317), .CLK(clk_in), .RSTB(n7286), .Q(
        \FIFO[101][18] ) );
  DFFARX1 \FIFO_reg[101][17]  ( .D(n1316), .CLK(clk_in), .RSTB(n7287), .Q(
        \FIFO[101][17] ) );
  DFFARX1 \FIFO_reg[101][16]  ( .D(n1315), .CLK(clk_in), .RSTB(n7287), .Q(
        \FIFO[101][16] ) );
  DFFARX1 \FIFO_reg[101][15]  ( .D(n1314), .CLK(clk_in), .RSTB(n7287), .Q(
        \FIFO[101][15] ) );
  DFFARX1 \FIFO_reg[101][14]  ( .D(n1313), .CLK(clk_in), .RSTB(n7287), .Q(
        \FIFO[101][14] ) );
  DFFARX1 \FIFO_reg[101][13]  ( .D(n1312), .CLK(clk_in), .RSTB(n7287), .Q(
        \FIFO[101][13] ) );
  DFFARX1 \FIFO_reg[101][12]  ( .D(n1311), .CLK(clk_in), .RSTB(n7287), .Q(
        \FIFO[101][12] ) );
  DFFARX1 \FIFO_reg[101][11]  ( .D(n1310), .CLK(clk_in), .RSTB(n7287), .Q(
        \FIFO[101][11] ) );
  DFFARX1 \FIFO_reg[101][10]  ( .D(n1309), .CLK(clk_in), .RSTB(n7287), .Q(
        \FIFO[101][10] ) );
  DFFARX1 \FIFO_reg[101][9]  ( .D(n1308), .CLK(clk_in), .RSTB(n7287), .Q(
        \FIFO[101][9] ) );
  DFFARX1 \FIFO_reg[101][8]  ( .D(n1307), .CLK(clk_in), .RSTB(n7287), .Q(
        \FIFO[101][8] ) );
  DFFARX1 \FIFO_reg[101][7]  ( .D(n1306), .CLK(clk_in), .RSTB(n7287), .Q(
        \FIFO[101][7] ) );
  DFFARX1 \FIFO_reg[101][6]  ( .D(n1305), .CLK(clk_in), .RSTB(n7287), .Q(
        \FIFO[101][6] ) );
  DFFARX1 \FIFO_reg[101][5]  ( .D(n1304), .CLK(clk_in), .RSTB(n7287), .Q(
        \FIFO[101][5] ) );
  DFFARX1 \FIFO_reg[101][4]  ( .D(n1303), .CLK(clk_in), .RSTB(n7287), .Q(
        \FIFO[101][4] ) );
  DFFARX1 \FIFO_reg[101][3]  ( .D(n1302), .CLK(clk_in), .RSTB(n7287), .Q(
        \FIFO[101][3] ) );
  DFFARX1 \FIFO_reg[101][2]  ( .D(n1301), .CLK(clk_in), .RSTB(n7287), .Q(
        \FIFO[101][2] ) );
  DFFARX1 \FIFO_reg[101][1]  ( .D(n1300), .CLK(clk_in), .RSTB(n7287), .Q(
        \FIFO[101][1] ) );
  DFFARX1 \FIFO_reg[101][0]  ( .D(n1299), .CLK(clk_in), .RSTB(n7287), .Q(
        \FIFO[101][0] ) );
  DFFARX1 \FIFO_reg[102][31]  ( .D(n1298), .CLK(clk_in), .RSTB(n7288), .Q(
        \FIFO[102][31] ) );
  DFFARX1 \FIFO_reg[102][30]  ( .D(n1297), .CLK(clk_in), .RSTB(n7288), .Q(
        \FIFO[102][30] ) );
  DFFARX1 \FIFO_reg[102][29]  ( .D(n1296), .CLK(clk_in), .RSTB(n7288), .Q(
        \FIFO[102][29] ) );
  DFFARX1 \FIFO_reg[102][28]  ( .D(n1295), .CLK(clk_in), .RSTB(n7288), .Q(
        \FIFO[102][28] ) );
  DFFARX1 \FIFO_reg[102][27]  ( .D(n1294), .CLK(clk_in), .RSTB(n7288), .Q(
        \FIFO[102][27] ) );
  DFFARX1 \FIFO_reg[102][26]  ( .D(n1293), .CLK(clk_in), .RSTB(n7288), .Q(
        \FIFO[102][26] ) );
  DFFARX1 \FIFO_reg[102][25]  ( .D(n1292), .CLK(clk_in), .RSTB(n7288), .Q(
        \FIFO[102][25] ) );
  DFFARX1 \FIFO_reg[102][24]  ( .D(n1291), .CLK(clk_in), .RSTB(n7288), .Q(
        \FIFO[102][24] ) );
  DFFARX1 \FIFO_reg[102][23]  ( .D(n1290), .CLK(clk_in), .RSTB(n7288), .Q(
        \FIFO[102][23] ) );
  DFFARX1 \FIFO_reg[102][22]  ( .D(n1289), .CLK(clk_in), .RSTB(n7288), .Q(
        \FIFO[102][22] ) );
  DFFARX1 \FIFO_reg[102][21]  ( .D(n1288), .CLK(clk_in), .RSTB(n7288), .Q(
        \FIFO[102][21] ) );
  DFFARX1 \FIFO_reg[102][20]  ( .D(n1287), .CLK(clk_in), .RSTB(n7288), .Q(
        \FIFO[102][20] ) );
  DFFARX1 \FIFO_reg[102][19]  ( .D(n1286), .CLK(clk_in), .RSTB(n7288), .Q(
        \FIFO[102][19] ) );
  DFFARX1 \FIFO_reg[102][18]  ( .D(n1285), .CLK(clk_in), .RSTB(n7288), .Q(
        \FIFO[102][18] ) );
  DFFARX1 \FIFO_reg[102][17]  ( .D(n1284), .CLK(clk_in), .RSTB(n7288), .Q(
        \FIFO[102][17] ) );
  DFFARX1 \FIFO_reg[102][16]  ( .D(n1283), .CLK(clk_in), .RSTB(n7288), .Q(
        \FIFO[102][16] ) );
  DFFARX1 \FIFO_reg[102][15]  ( .D(n1282), .CLK(clk_in), .RSTB(n7288), .Q(
        \FIFO[102][15] ) );
  DFFARX1 \FIFO_reg[102][14]  ( .D(n1281), .CLK(clk_in), .RSTB(n7288), .Q(
        \FIFO[102][14] ) );
  DFFARX1 \FIFO_reg[102][13]  ( .D(n1280), .CLK(clk_in), .RSTB(n7289), .Q(
        \FIFO[102][13] ) );
  DFFARX1 \FIFO_reg[102][12]  ( .D(n1279), .CLK(clk_in), .RSTB(n7289), .Q(
        \FIFO[102][12] ) );
  DFFARX1 \FIFO_reg[102][11]  ( .D(n1278), .CLK(clk_in), .RSTB(n7289), .Q(
        \FIFO[102][11] ) );
  DFFARX1 \FIFO_reg[102][10]  ( .D(n1277), .CLK(clk_in), .RSTB(n7289), .Q(
        \FIFO[102][10] ) );
  DFFARX1 \FIFO_reg[102][9]  ( .D(n1276), .CLK(clk_in), .RSTB(n7289), .Q(
        \FIFO[102][9] ) );
  DFFARX1 \FIFO_reg[102][8]  ( .D(n1275), .CLK(clk_in), .RSTB(n7289), .Q(
        \FIFO[102][8] ) );
  DFFARX1 \FIFO_reg[102][7]  ( .D(n1274), .CLK(clk_in), .RSTB(n7289), .Q(
        \FIFO[102][7] ) );
  DFFARX1 \FIFO_reg[102][6]  ( .D(n1273), .CLK(clk_in), .RSTB(n7289), .Q(
        \FIFO[102][6] ) );
  DFFARX1 \FIFO_reg[102][5]  ( .D(n1272), .CLK(clk_in), .RSTB(n7289), .Q(
        \FIFO[102][5] ) );
  DFFARX1 \FIFO_reg[102][4]  ( .D(n1271), .CLK(clk_in), .RSTB(n7289), .Q(
        \FIFO[102][4] ) );
  DFFARX1 \FIFO_reg[102][3]  ( .D(n1270), .CLK(clk_in), .RSTB(n7289), .Q(
        \FIFO[102][3] ) );
  DFFARX1 \FIFO_reg[102][2]  ( .D(n1269), .CLK(clk_in), .RSTB(n7289), .Q(
        \FIFO[102][2] ) );
  DFFARX1 \FIFO_reg[102][1]  ( .D(n1268), .CLK(clk_in), .RSTB(n7289), .Q(
        \FIFO[102][1] ) );
  DFFARX1 \FIFO_reg[102][0]  ( .D(n1267), .CLK(clk_in), .RSTB(n7289), .Q(
        \FIFO[102][0] ) );
  DFFARX1 \FIFO_reg[103][31]  ( .D(n1266), .CLK(clk_in), .RSTB(n7289), .Q(
        \FIFO[103][31] ) );
  DFFARX1 \FIFO_reg[103][30]  ( .D(n1265), .CLK(clk_in), .RSTB(n7289), .Q(
        \FIFO[103][30] ) );
  DFFARX1 \FIFO_reg[103][29]  ( .D(n1264), .CLK(clk_in), .RSTB(n7289), .Q(
        \FIFO[103][29] ) );
  DFFARX1 \FIFO_reg[103][28]  ( .D(n1263), .CLK(clk_in), .RSTB(n7289), .Q(
        \FIFO[103][28] ) );
  DFFARX1 \FIFO_reg[103][27]  ( .D(n1262), .CLK(clk_in), .RSTB(n7290), .Q(
        \FIFO[103][27] ) );
  DFFARX1 \FIFO_reg[103][26]  ( .D(n1261), .CLK(clk_in), .RSTB(n7290), .Q(
        \FIFO[103][26] ) );
  DFFARX1 \FIFO_reg[103][25]  ( .D(n1260), .CLK(clk_in), .RSTB(n7290), .Q(
        \FIFO[103][25] ) );
  DFFARX1 \FIFO_reg[103][24]  ( .D(n1259), .CLK(clk_in), .RSTB(n7290), .Q(
        \FIFO[103][24] ) );
  DFFARX1 \FIFO_reg[103][23]  ( .D(n1258), .CLK(clk_in), .RSTB(n7290), .Q(
        \FIFO[103][23] ) );
  DFFARX1 \FIFO_reg[103][22]  ( .D(n1257), .CLK(clk_in), .RSTB(n7290), .Q(
        \FIFO[103][22] ) );
  DFFARX1 \FIFO_reg[103][21]  ( .D(n1256), .CLK(clk_in), .RSTB(n7290), .Q(
        \FIFO[103][21] ) );
  DFFARX1 \FIFO_reg[103][20]  ( .D(n1255), .CLK(clk_in), .RSTB(n7290), .Q(
        \FIFO[103][20] ) );
  DFFARX1 \FIFO_reg[103][19]  ( .D(n1254), .CLK(clk_in), .RSTB(n7290), .Q(
        \FIFO[103][19] ) );
  DFFARX1 \FIFO_reg[103][18]  ( .D(n1253), .CLK(clk_in), .RSTB(n7290), .Q(
        \FIFO[103][18] ) );
  DFFARX1 \FIFO_reg[103][17]  ( .D(n1252), .CLK(clk_in), .RSTB(n7290), .Q(
        \FIFO[103][17] ) );
  DFFARX1 \FIFO_reg[103][16]  ( .D(n1251), .CLK(clk_in), .RSTB(n7290), .Q(
        \FIFO[103][16] ) );
  DFFARX1 \FIFO_reg[103][15]  ( .D(n1250), .CLK(clk_in), .RSTB(n7290), .Q(
        \FIFO[103][15] ) );
  DFFARX1 \FIFO_reg[103][14]  ( .D(n1249), .CLK(clk_in), .RSTB(n7290), .Q(
        \FIFO[103][14] ) );
  DFFARX1 \FIFO_reg[103][13]  ( .D(n1248), .CLK(clk_in), .RSTB(n7290), .Q(
        \FIFO[103][13] ) );
  DFFARX1 \FIFO_reg[103][12]  ( .D(n1247), .CLK(clk_in), .RSTB(n7290), .Q(
        \FIFO[103][12] ) );
  DFFARX1 \FIFO_reg[103][11]  ( .D(n1246), .CLK(clk_in), .RSTB(n7290), .Q(
        \FIFO[103][11] ) );
  DFFARX1 \FIFO_reg[103][10]  ( .D(n1245), .CLK(clk_in), .RSTB(n7290), .Q(
        \FIFO[103][10] ) );
  DFFARX1 \FIFO_reg[103][9]  ( .D(n1244), .CLK(clk_in), .RSTB(n7291), .Q(
        \FIFO[103][9] ) );
  DFFARX1 \FIFO_reg[103][8]  ( .D(n1243), .CLK(clk_in), .RSTB(n7291), .Q(
        \FIFO[103][8] ) );
  DFFARX1 \FIFO_reg[103][7]  ( .D(n1242), .CLK(clk_in), .RSTB(n7291), .Q(
        \FIFO[103][7] ) );
  DFFARX1 \FIFO_reg[103][6]  ( .D(n1241), .CLK(clk_in), .RSTB(n7291), .Q(
        \FIFO[103][6] ) );
  DFFARX1 \FIFO_reg[103][5]  ( .D(n1240), .CLK(clk_in), .RSTB(n7291), .Q(
        \FIFO[103][5] ) );
  DFFARX1 \FIFO_reg[103][4]  ( .D(n1239), .CLK(clk_in), .RSTB(n7291), .Q(
        \FIFO[103][4] ) );
  DFFARX1 \FIFO_reg[103][3]  ( .D(n1238), .CLK(clk_in), .RSTB(n7291), .Q(
        \FIFO[103][3] ) );
  DFFARX1 \FIFO_reg[103][2]  ( .D(n1237), .CLK(clk_in), .RSTB(n7291), .Q(
        \FIFO[103][2] ) );
  DFFARX1 \FIFO_reg[103][1]  ( .D(n1236), .CLK(clk_in), .RSTB(n7291), .Q(
        \FIFO[103][1] ) );
  DFFARX1 \FIFO_reg[103][0]  ( .D(n1235), .CLK(clk_in), .RSTB(n7291), .Q(
        \FIFO[103][0] ) );
  DFFARX1 \FIFO_reg[104][31]  ( .D(n1234), .CLK(clk_in), .RSTB(n7291), .Q(
        \FIFO[104][31] ) );
  DFFARX1 \FIFO_reg[104][30]  ( .D(n1233), .CLK(clk_in), .RSTB(n7291), .Q(
        \FIFO[104][30] ) );
  DFFARX1 \FIFO_reg[104][29]  ( .D(n1232), .CLK(clk_in), .RSTB(n7291), .Q(
        \FIFO[104][29] ) );
  DFFARX1 \FIFO_reg[104][28]  ( .D(n1231), .CLK(clk_in), .RSTB(n7291), .Q(
        \FIFO[104][28] ) );
  DFFARX1 \FIFO_reg[104][27]  ( .D(n1230), .CLK(clk_in), .RSTB(n7291), .Q(
        \FIFO[104][27] ) );
  DFFARX1 \FIFO_reg[104][26]  ( .D(n1229), .CLK(clk_in), .RSTB(n7291), .Q(
        \FIFO[104][26] ) );
  DFFARX1 \FIFO_reg[104][25]  ( .D(n1228), .CLK(clk_in), .RSTB(n7291), .Q(
        \FIFO[104][25] ) );
  DFFARX1 \FIFO_reg[104][24]  ( .D(n1227), .CLK(clk_in), .RSTB(n7291), .Q(
        \FIFO[104][24] ) );
  DFFARX1 \FIFO_reg[104][23]  ( .D(n1226), .CLK(clk_in), .RSTB(n7292), .Q(
        \FIFO[104][23] ) );
  DFFARX1 \FIFO_reg[104][22]  ( .D(n1225), .CLK(clk_in), .RSTB(n7292), .Q(
        \FIFO[104][22] ) );
  DFFARX1 \FIFO_reg[104][21]  ( .D(n1224), .CLK(clk_in), .RSTB(n7292), .Q(
        \FIFO[104][21] ) );
  DFFARX1 \FIFO_reg[104][20]  ( .D(n1223), .CLK(clk_in), .RSTB(n7292), .Q(
        \FIFO[104][20] ) );
  DFFARX1 \FIFO_reg[104][19]  ( .D(n1222), .CLK(clk_in), .RSTB(n7292), .Q(
        \FIFO[104][19] ) );
  DFFARX1 \FIFO_reg[104][18]  ( .D(n1221), .CLK(clk_in), .RSTB(n7292), .Q(
        \FIFO[104][18] ) );
  DFFARX1 \FIFO_reg[104][17]  ( .D(n1220), .CLK(clk_in), .RSTB(n7292), .Q(
        \FIFO[104][17] ) );
  DFFARX1 \FIFO_reg[104][16]  ( .D(n1219), .CLK(clk_in), .RSTB(n7292), .Q(
        \FIFO[104][16] ) );
  DFFARX1 \FIFO_reg[104][15]  ( .D(n1218), .CLK(clk_in), .RSTB(n7292), .Q(
        \FIFO[104][15] ) );
  DFFARX1 \FIFO_reg[104][14]  ( .D(n1217), .CLK(clk_in), .RSTB(n7292), .Q(
        \FIFO[104][14] ) );
  DFFARX1 \FIFO_reg[104][13]  ( .D(n1216), .CLK(clk_in), .RSTB(n7292), .Q(
        \FIFO[104][13] ) );
  DFFARX1 \FIFO_reg[104][12]  ( .D(n1215), .CLK(clk_in), .RSTB(n7292), .Q(
        \FIFO[104][12] ) );
  DFFARX1 \FIFO_reg[104][11]  ( .D(n1214), .CLK(clk_in), .RSTB(n7292), .Q(
        \FIFO[104][11] ) );
  DFFARX1 \FIFO_reg[104][10]  ( .D(n1213), .CLK(clk_in), .RSTB(n7292), .Q(
        \FIFO[104][10] ) );
  DFFARX1 \FIFO_reg[104][9]  ( .D(n1212), .CLK(clk_in), .RSTB(n7292), .Q(
        \FIFO[104][9] ) );
  DFFARX1 \FIFO_reg[104][8]  ( .D(n1211), .CLK(clk_in), .RSTB(n7292), .Q(
        \FIFO[104][8] ) );
  DFFARX1 \FIFO_reg[104][7]  ( .D(n1210), .CLK(clk_in), .RSTB(n7292), .Q(
        \FIFO[104][7] ) );
  DFFARX1 \FIFO_reg[104][6]  ( .D(n1209), .CLK(clk_in), .RSTB(n7292), .Q(
        \FIFO[104][6] ) );
  DFFARX1 \FIFO_reg[104][5]  ( .D(n1208), .CLK(clk_in), .RSTB(n7293), .Q(
        \FIFO[104][5] ) );
  DFFARX1 \FIFO_reg[104][4]  ( .D(n1207), .CLK(clk_in), .RSTB(n7293), .Q(
        \FIFO[104][4] ) );
  DFFARX1 \FIFO_reg[104][3]  ( .D(n1206), .CLK(clk_in), .RSTB(n7293), .Q(
        \FIFO[104][3] ) );
  DFFARX1 \FIFO_reg[104][2]  ( .D(n1205), .CLK(clk_in), .RSTB(n7293), .Q(
        \FIFO[104][2] ) );
  DFFARX1 \FIFO_reg[104][1]  ( .D(n1204), .CLK(clk_in), .RSTB(n7293), .Q(
        \FIFO[104][1] ) );
  DFFARX1 \FIFO_reg[104][0]  ( .D(n1203), .CLK(clk_in), .RSTB(n7293), .Q(
        \FIFO[104][0] ) );
  DFFARX1 \FIFO_reg[105][31]  ( .D(n1202), .CLK(clk_in), .RSTB(n7293), .Q(
        \FIFO[105][31] ) );
  DFFARX1 \FIFO_reg[105][30]  ( .D(n1201), .CLK(clk_in), .RSTB(n7293), .Q(
        \FIFO[105][30] ) );
  DFFARX1 \FIFO_reg[105][29]  ( .D(n1200), .CLK(clk_in), .RSTB(n7293), .Q(
        \FIFO[105][29] ) );
  DFFARX1 \FIFO_reg[105][28]  ( .D(n1199), .CLK(clk_in), .RSTB(n7293), .Q(
        \FIFO[105][28] ) );
  DFFARX1 \FIFO_reg[105][27]  ( .D(n1198), .CLK(clk_in), .RSTB(n7293), .Q(
        \FIFO[105][27] ) );
  DFFARX1 \FIFO_reg[105][26]  ( .D(n1197), .CLK(clk_in), .RSTB(n7293), .Q(
        \FIFO[105][26] ) );
  DFFARX1 \FIFO_reg[105][25]  ( .D(n1196), .CLK(clk_in), .RSTB(n7293), .Q(
        \FIFO[105][25] ) );
  DFFARX1 \FIFO_reg[105][24]  ( .D(n1195), .CLK(clk_in), .RSTB(n7293), .Q(
        \FIFO[105][24] ) );
  DFFARX1 \FIFO_reg[105][23]  ( .D(n1194), .CLK(clk_in), .RSTB(n7293), .Q(
        \FIFO[105][23] ) );
  DFFARX1 \FIFO_reg[105][22]  ( .D(n1193), .CLK(clk_in), .RSTB(n7293), .Q(
        \FIFO[105][22] ) );
  DFFARX1 \FIFO_reg[105][21]  ( .D(n1192), .CLK(clk_in), .RSTB(n7293), .Q(
        \FIFO[105][21] ) );
  DFFARX1 \FIFO_reg[105][20]  ( .D(n1191), .CLK(clk_in), .RSTB(n7293), .Q(
        \FIFO[105][20] ) );
  DFFARX1 \FIFO_reg[105][19]  ( .D(n1190), .CLK(clk_in), .RSTB(n7294), .Q(
        \FIFO[105][19] ) );
  DFFARX1 \FIFO_reg[105][18]  ( .D(n1189), .CLK(clk_in), .RSTB(n7294), .Q(
        \FIFO[105][18] ) );
  DFFARX1 \FIFO_reg[105][17]  ( .D(n1188), .CLK(clk_in), .RSTB(n7294), .Q(
        \FIFO[105][17] ) );
  DFFARX1 \FIFO_reg[105][16]  ( .D(n1187), .CLK(clk_in), .RSTB(n7294), .Q(
        \FIFO[105][16] ) );
  DFFARX1 \FIFO_reg[105][15]  ( .D(n1186), .CLK(clk_in), .RSTB(n7294), .Q(
        \FIFO[105][15] ) );
  DFFARX1 \FIFO_reg[105][14]  ( .D(n1185), .CLK(clk_in), .RSTB(n7294), .Q(
        \FIFO[105][14] ) );
  DFFARX1 \FIFO_reg[105][13]  ( .D(n1184), .CLK(clk_in), .RSTB(n7294), .Q(
        \FIFO[105][13] ) );
  DFFARX1 \FIFO_reg[105][12]  ( .D(n1183), .CLK(clk_in), .RSTB(n7294), .Q(
        \FIFO[105][12] ) );
  DFFARX1 \FIFO_reg[105][11]  ( .D(n1182), .CLK(clk_in), .RSTB(n7294), .Q(
        \FIFO[105][11] ) );
  DFFARX1 \FIFO_reg[105][10]  ( .D(n1181), .CLK(clk_in), .RSTB(n7294), .Q(
        \FIFO[105][10] ) );
  DFFARX1 \FIFO_reg[105][9]  ( .D(n1180), .CLK(clk_in), .RSTB(n7294), .Q(
        \FIFO[105][9] ) );
  DFFARX1 \FIFO_reg[105][8]  ( .D(n1179), .CLK(clk_in), .RSTB(n7294), .Q(
        \FIFO[105][8] ) );
  DFFARX1 \FIFO_reg[105][7]  ( .D(n1178), .CLK(clk_in), .RSTB(n7294), .Q(
        \FIFO[105][7] ) );
  DFFARX1 \FIFO_reg[105][6]  ( .D(n1177), .CLK(clk_in), .RSTB(n7294), .Q(
        \FIFO[105][6] ) );
  DFFARX1 \FIFO_reg[105][5]  ( .D(n1176), .CLK(clk_in), .RSTB(n7294), .Q(
        \FIFO[105][5] ) );
  DFFARX1 \FIFO_reg[105][4]  ( .D(n1175), .CLK(clk_in), .RSTB(n7294), .Q(
        \FIFO[105][4] ) );
  DFFARX1 \FIFO_reg[105][3]  ( .D(n1174), .CLK(clk_in), .RSTB(n7294), .Q(
        \FIFO[105][3] ) );
  DFFARX1 \FIFO_reg[105][2]  ( .D(n1173), .CLK(clk_in), .RSTB(n7294), .Q(
        \FIFO[105][2] ) );
  DFFARX1 \FIFO_reg[105][1]  ( .D(n1172), .CLK(clk_in), .RSTB(n7295), .Q(
        \FIFO[105][1] ) );
  DFFARX1 \FIFO_reg[105][0]  ( .D(n1171), .CLK(clk_in), .RSTB(n7295), .Q(
        \FIFO[105][0] ) );
  DFFARX1 \FIFO_reg[106][31]  ( .D(n1170), .CLK(clk_in), .RSTB(n7295), .Q(
        \FIFO[106][31] ) );
  DFFARX1 \FIFO_reg[106][30]  ( .D(n1169), .CLK(clk_in), .RSTB(n7295), .Q(
        \FIFO[106][30] ) );
  DFFARX1 \FIFO_reg[106][29]  ( .D(n1168), .CLK(clk_in), .RSTB(n7295), .Q(
        \FIFO[106][29] ) );
  DFFARX1 \FIFO_reg[106][28]  ( .D(n1167), .CLK(clk_in), .RSTB(n7295), .Q(
        \FIFO[106][28] ) );
  DFFARX1 \FIFO_reg[106][27]  ( .D(n1166), .CLK(clk_in), .RSTB(n7295), .Q(
        \FIFO[106][27] ) );
  DFFARX1 \FIFO_reg[106][26]  ( .D(n1165), .CLK(clk_in), .RSTB(n7295), .Q(
        \FIFO[106][26] ) );
  DFFARX1 \FIFO_reg[106][25]  ( .D(n1164), .CLK(clk_in), .RSTB(n7295), .Q(
        \FIFO[106][25] ) );
  DFFARX1 \FIFO_reg[106][24]  ( .D(n1163), .CLK(clk_in), .RSTB(n7295), .Q(
        \FIFO[106][24] ) );
  DFFARX1 \FIFO_reg[106][23]  ( .D(n1162), .CLK(clk_in), .RSTB(n7295), .Q(
        \FIFO[106][23] ) );
  DFFARX1 \FIFO_reg[106][22]  ( .D(n1161), .CLK(clk_in), .RSTB(n7295), .Q(
        \FIFO[106][22] ) );
  DFFARX1 \FIFO_reg[106][21]  ( .D(n1160), .CLK(clk_in), .RSTB(n7295), .Q(
        \FIFO[106][21] ) );
  DFFARX1 \FIFO_reg[106][20]  ( .D(n1159), .CLK(clk_in), .RSTB(n7295), .Q(
        \FIFO[106][20] ) );
  DFFARX1 \FIFO_reg[106][19]  ( .D(n1158), .CLK(clk_in), .RSTB(n7295), .Q(
        \FIFO[106][19] ) );
  DFFARX1 \FIFO_reg[106][18]  ( .D(n1157), .CLK(clk_in), .RSTB(n7295), .Q(
        \FIFO[106][18] ) );
  DFFARX1 \FIFO_reg[106][17]  ( .D(n1156), .CLK(clk_in), .RSTB(n7295), .Q(
        \FIFO[106][17] ) );
  DFFARX1 \FIFO_reg[106][16]  ( .D(n1155), .CLK(clk_in), .RSTB(n7295), .Q(
        \FIFO[106][16] ) );
  DFFARX1 \FIFO_reg[106][15]  ( .D(n1154), .CLK(clk_in), .RSTB(n7296), .Q(
        \FIFO[106][15] ) );
  DFFARX1 \FIFO_reg[106][14]  ( .D(n1153), .CLK(clk_in), .RSTB(n7296), .Q(
        \FIFO[106][14] ) );
  DFFARX1 \FIFO_reg[106][13]  ( .D(n1152), .CLK(clk_in), .RSTB(n7296), .Q(
        \FIFO[106][13] ) );
  DFFARX1 \FIFO_reg[106][12]  ( .D(n1151), .CLK(clk_in), .RSTB(n7296), .Q(
        \FIFO[106][12] ) );
  DFFARX1 \FIFO_reg[106][11]  ( .D(n1150), .CLK(clk_in), .RSTB(n7296), .Q(
        \FIFO[106][11] ) );
  DFFARX1 \FIFO_reg[106][10]  ( .D(n1149), .CLK(clk_in), .RSTB(n7296), .Q(
        \FIFO[106][10] ) );
  DFFARX1 \FIFO_reg[106][9]  ( .D(n1148), .CLK(clk_in), .RSTB(n7296), .Q(
        \FIFO[106][9] ) );
  DFFARX1 \FIFO_reg[106][8]  ( .D(n1147), .CLK(clk_in), .RSTB(n7296), .Q(
        \FIFO[106][8] ) );
  DFFARX1 \FIFO_reg[106][7]  ( .D(n1146), .CLK(clk_in), .RSTB(n7296), .Q(
        \FIFO[106][7] ) );
  DFFARX1 \FIFO_reg[106][6]  ( .D(n1145), .CLK(clk_in), .RSTB(n7296), .Q(
        \FIFO[106][6] ) );
  DFFARX1 \FIFO_reg[106][5]  ( .D(n1144), .CLK(clk_in), .RSTB(n7296), .Q(
        \FIFO[106][5] ) );
  DFFARX1 \FIFO_reg[106][4]  ( .D(n1143), .CLK(clk_in), .RSTB(n7296), .Q(
        \FIFO[106][4] ) );
  DFFARX1 \FIFO_reg[106][3]  ( .D(n1142), .CLK(clk_in), .RSTB(n7296), .Q(
        \FIFO[106][3] ) );
  DFFARX1 \FIFO_reg[106][2]  ( .D(n1141), .CLK(clk_in), .RSTB(n7296), .Q(
        \FIFO[106][2] ) );
  DFFARX1 \FIFO_reg[106][1]  ( .D(n1140), .CLK(clk_in), .RSTB(n7296), .Q(
        \FIFO[106][1] ) );
  DFFARX1 \FIFO_reg[106][0]  ( .D(n1139), .CLK(clk_in), .RSTB(n7296), .Q(
        \FIFO[106][0] ) );
  DFFARX1 \FIFO_reg[107][31]  ( .D(n1138), .CLK(clk_in), .RSTB(n7296), .Q(
        \FIFO[107][31] ) );
  DFFARX1 \FIFO_reg[107][30]  ( .D(n1137), .CLK(clk_in), .RSTB(n7296), .Q(
        \FIFO[107][30] ) );
  DFFARX1 \FIFO_reg[107][29]  ( .D(n1136), .CLK(clk_in), .RSTB(n7297), .Q(
        \FIFO[107][29] ) );
  DFFARX1 \FIFO_reg[107][28]  ( .D(n1135), .CLK(clk_in), .RSTB(n7297), .Q(
        \FIFO[107][28] ) );
  DFFARX1 \FIFO_reg[107][27]  ( .D(n1134), .CLK(clk_in), .RSTB(n7297), .Q(
        \FIFO[107][27] ) );
  DFFARX1 \FIFO_reg[107][26]  ( .D(n1133), .CLK(clk_in), .RSTB(n7297), .Q(
        \FIFO[107][26] ) );
  DFFARX1 \FIFO_reg[107][25]  ( .D(n1132), .CLK(clk_in), .RSTB(n7297), .Q(
        \FIFO[107][25] ) );
  DFFARX1 \FIFO_reg[107][24]  ( .D(n1131), .CLK(clk_in), .RSTB(n7297), .Q(
        \FIFO[107][24] ) );
  DFFARX1 \FIFO_reg[107][23]  ( .D(n1130), .CLK(clk_in), .RSTB(n7297), .Q(
        \FIFO[107][23] ) );
  DFFARX1 \FIFO_reg[107][22]  ( .D(n1129), .CLK(clk_in), .RSTB(n7297), .Q(
        \FIFO[107][22] ) );
  DFFARX1 \FIFO_reg[107][21]  ( .D(n1128), .CLK(clk_in), .RSTB(n7297), .Q(
        \FIFO[107][21] ) );
  DFFARX1 \FIFO_reg[107][20]  ( .D(n1127), .CLK(clk_in), .RSTB(n7297), .Q(
        \FIFO[107][20] ) );
  DFFARX1 \FIFO_reg[107][19]  ( .D(n1126), .CLK(clk_in), .RSTB(n7297), .Q(
        \FIFO[107][19] ) );
  DFFARX1 \FIFO_reg[107][18]  ( .D(n1125), .CLK(clk_in), .RSTB(n7297), .Q(
        \FIFO[107][18] ) );
  DFFARX1 \FIFO_reg[107][17]  ( .D(n1124), .CLK(clk_in), .RSTB(n7297), .Q(
        \FIFO[107][17] ) );
  DFFARX1 \FIFO_reg[107][16]  ( .D(n1123), .CLK(clk_in), .RSTB(n7297), .Q(
        \FIFO[107][16] ) );
  DFFARX1 \FIFO_reg[107][15]  ( .D(n1122), .CLK(clk_in), .RSTB(n7297), .Q(
        \FIFO[107][15] ) );
  DFFARX1 \FIFO_reg[107][14]  ( .D(n1121), .CLK(clk_in), .RSTB(n7297), .Q(
        \FIFO[107][14] ) );
  DFFARX1 \FIFO_reg[107][13]  ( .D(n1120), .CLK(clk_in), .RSTB(n7297), .Q(
        \FIFO[107][13] ) );
  DFFARX1 \FIFO_reg[107][12]  ( .D(n1119), .CLK(clk_in), .RSTB(n7297), .Q(
        \FIFO[107][12] ) );
  DFFARX1 \FIFO_reg[107][11]  ( .D(n1118), .CLK(clk_in), .RSTB(n7298), .Q(
        \FIFO[107][11] ) );
  DFFARX1 \FIFO_reg[107][10]  ( .D(n1117), .CLK(clk_in), .RSTB(n7298), .Q(
        \FIFO[107][10] ) );
  DFFARX1 \FIFO_reg[107][9]  ( .D(n1116), .CLK(clk_in), .RSTB(n7298), .Q(
        \FIFO[107][9] ) );
  DFFARX1 \FIFO_reg[107][8]  ( .D(n1115), .CLK(clk_in), .RSTB(n7298), .Q(
        \FIFO[107][8] ) );
  DFFARX1 \FIFO_reg[107][7]  ( .D(n1114), .CLK(clk_in), .RSTB(n7298), .Q(
        \FIFO[107][7] ) );
  DFFARX1 \FIFO_reg[107][6]  ( .D(n1113), .CLK(clk_in), .RSTB(n7298), .Q(
        \FIFO[107][6] ) );
  DFFARX1 \FIFO_reg[107][5]  ( .D(n1112), .CLK(clk_in), .RSTB(n7298), .Q(
        \FIFO[107][5] ) );
  DFFARX1 \FIFO_reg[107][4]  ( .D(n1111), .CLK(clk_in), .RSTB(n7298), .Q(
        \FIFO[107][4] ) );
  DFFARX1 \FIFO_reg[107][3]  ( .D(n1110), .CLK(clk_in), .RSTB(n7298), .Q(
        \FIFO[107][3] ) );
  DFFARX1 \FIFO_reg[107][2]  ( .D(n1109), .CLK(clk_in), .RSTB(n7298), .Q(
        \FIFO[107][2] ) );
  DFFARX1 \FIFO_reg[107][1]  ( .D(n1108), .CLK(clk_in), .RSTB(n7298), .Q(
        \FIFO[107][1] ) );
  DFFARX1 \FIFO_reg[107][0]  ( .D(n1107), .CLK(clk_in), .RSTB(n7298), .Q(
        \FIFO[107][0] ) );
  DFFARX1 \FIFO_reg[108][31]  ( .D(n1106), .CLK(clk_in), .RSTB(n7298), .Q(
        \FIFO[108][31] ) );
  DFFARX1 \FIFO_reg[108][30]  ( .D(n1105), .CLK(clk_in), .RSTB(n7298), .Q(
        \FIFO[108][30] ) );
  DFFARX1 \FIFO_reg[108][29]  ( .D(n1104), .CLK(clk_in), .RSTB(n7298), .Q(
        \FIFO[108][29] ) );
  DFFARX1 \FIFO_reg[108][28]  ( .D(n1103), .CLK(clk_in), .RSTB(n7298), .Q(
        \FIFO[108][28] ) );
  DFFARX1 \FIFO_reg[108][27]  ( .D(n1102), .CLK(clk_in), .RSTB(n7298), .Q(
        \FIFO[108][27] ) );
  DFFARX1 \FIFO_reg[108][26]  ( .D(n1101), .CLK(clk_in), .RSTB(n7298), .Q(
        \FIFO[108][26] ) );
  DFFARX1 \FIFO_reg[108][25]  ( .D(n1100), .CLK(clk_in), .RSTB(n7299), .Q(
        \FIFO[108][25] ) );
  DFFARX1 \FIFO_reg[108][24]  ( .D(n1099), .CLK(clk_in), .RSTB(n7299), .Q(
        \FIFO[108][24] ) );
  DFFARX1 \FIFO_reg[108][23]  ( .D(n1098), .CLK(clk_in), .RSTB(n7299), .Q(
        \FIFO[108][23] ) );
  DFFARX1 \FIFO_reg[108][22]  ( .D(n1097), .CLK(clk_in), .RSTB(n7299), .Q(
        \FIFO[108][22] ) );
  DFFARX1 \FIFO_reg[108][21]  ( .D(n1096), .CLK(clk_in), .RSTB(n7299), .Q(
        \FIFO[108][21] ) );
  DFFARX1 \FIFO_reg[108][20]  ( .D(n1095), .CLK(clk_in), .RSTB(n7299), .Q(
        \FIFO[108][20] ) );
  DFFARX1 \FIFO_reg[108][19]  ( .D(n1094), .CLK(clk_in), .RSTB(n7299), .Q(
        \FIFO[108][19] ) );
  DFFARX1 \FIFO_reg[108][18]  ( .D(n1093), .CLK(clk_in), .RSTB(n7299), .Q(
        \FIFO[108][18] ) );
  DFFARX1 \FIFO_reg[108][17]  ( .D(n1092), .CLK(clk_in), .RSTB(n7299), .Q(
        \FIFO[108][17] ) );
  DFFARX1 \FIFO_reg[108][16]  ( .D(n1091), .CLK(clk_in), .RSTB(n7299), .Q(
        \FIFO[108][16] ) );
  DFFARX1 \FIFO_reg[108][15]  ( .D(n1090), .CLK(clk_in), .RSTB(n7299), .Q(
        \FIFO[108][15] ) );
  DFFARX1 \FIFO_reg[108][14]  ( .D(n1089), .CLK(clk_in), .RSTB(n7299), .Q(
        \FIFO[108][14] ) );
  DFFARX1 \FIFO_reg[108][13]  ( .D(n1088), .CLK(clk_in), .RSTB(n7299), .Q(
        \FIFO[108][13] ) );
  DFFARX1 \FIFO_reg[108][12]  ( .D(n1087), .CLK(clk_in), .RSTB(n7299), .Q(
        \FIFO[108][12] ) );
  DFFARX1 \FIFO_reg[108][11]  ( .D(n1086), .CLK(clk_in), .RSTB(n7299), .Q(
        \FIFO[108][11] ) );
  DFFARX1 \FIFO_reg[108][10]  ( .D(n1085), .CLK(clk_in), .RSTB(n7299), .Q(
        \FIFO[108][10] ) );
  DFFARX1 \FIFO_reg[108][9]  ( .D(n1084), .CLK(clk_in), .RSTB(n7299), .Q(
        \FIFO[108][9] ) );
  DFFARX1 \FIFO_reg[108][8]  ( .D(n1083), .CLK(clk_in), .RSTB(n7299), .Q(
        \FIFO[108][8] ) );
  DFFARX1 \FIFO_reg[108][7]  ( .D(n1082), .CLK(clk_in), .RSTB(n7300), .Q(
        \FIFO[108][7] ) );
  DFFARX1 \FIFO_reg[108][6]  ( .D(n1081), .CLK(clk_in), .RSTB(n7300), .Q(
        \FIFO[108][6] ) );
  DFFARX1 \FIFO_reg[108][5]  ( .D(n1080), .CLK(clk_in), .RSTB(n7300), .Q(
        \FIFO[108][5] ) );
  DFFARX1 \FIFO_reg[108][4]  ( .D(n1079), .CLK(clk_in), .RSTB(n7300), .Q(
        \FIFO[108][4] ) );
  DFFARX1 \FIFO_reg[108][3]  ( .D(n1078), .CLK(clk_in), .RSTB(n7300), .Q(
        \FIFO[108][3] ) );
  DFFARX1 \FIFO_reg[108][2]  ( .D(n1077), .CLK(clk_in), .RSTB(n7300), .Q(
        \FIFO[108][2] ) );
  DFFARX1 \FIFO_reg[108][1]  ( .D(n1076), .CLK(clk_in), .RSTB(n7300), .Q(
        \FIFO[108][1] ) );
  DFFARX1 \FIFO_reg[108][0]  ( .D(n1075), .CLK(clk_in), .RSTB(n7300), .Q(
        \FIFO[108][0] ) );
  DFFARX1 \FIFO_reg[109][31]  ( .D(n1074), .CLK(clk_in), .RSTB(n7300), .Q(
        \FIFO[109][31] ) );
  DFFARX1 \FIFO_reg[109][30]  ( .D(n1073), .CLK(clk_in), .RSTB(n7300), .Q(
        \FIFO[109][30] ) );
  DFFARX1 \FIFO_reg[109][29]  ( .D(n1072), .CLK(clk_in), .RSTB(n7300), .Q(
        \FIFO[109][29] ) );
  DFFARX1 \FIFO_reg[109][28]  ( .D(n1071), .CLK(clk_in), .RSTB(n7300), .Q(
        \FIFO[109][28] ) );
  DFFARX1 \FIFO_reg[109][27]  ( .D(n1070), .CLK(clk_in), .RSTB(n7300), .Q(
        \FIFO[109][27] ) );
  DFFARX1 \FIFO_reg[109][26]  ( .D(n1069), .CLK(clk_in), .RSTB(n7300), .Q(
        \FIFO[109][26] ) );
  DFFARX1 \FIFO_reg[109][25]  ( .D(n1068), .CLK(clk_in), .RSTB(n7300), .Q(
        \FIFO[109][25] ) );
  DFFARX1 \FIFO_reg[109][24]  ( .D(n1067), .CLK(clk_in), .RSTB(n7300), .Q(
        \FIFO[109][24] ) );
  DFFARX1 \FIFO_reg[109][23]  ( .D(n1066), .CLK(clk_in), .RSTB(n7300), .Q(
        \FIFO[109][23] ) );
  DFFARX1 \FIFO_reg[109][22]  ( .D(n1065), .CLK(clk_in), .RSTB(n7300), .Q(
        \FIFO[109][22] ) );
  DFFARX1 \FIFO_reg[109][21]  ( .D(n1064), .CLK(clk_in), .RSTB(n7301), .Q(
        \FIFO[109][21] ) );
  DFFARX1 \FIFO_reg[109][20]  ( .D(n1063), .CLK(clk_in), .RSTB(n7301), .Q(
        \FIFO[109][20] ) );
  DFFARX1 \FIFO_reg[109][19]  ( .D(n1062), .CLK(clk_in), .RSTB(n7301), .Q(
        \FIFO[109][19] ) );
  DFFARX1 \FIFO_reg[109][18]  ( .D(n1061), .CLK(clk_in), .RSTB(n7301), .Q(
        \FIFO[109][18] ) );
  DFFARX1 \FIFO_reg[109][17]  ( .D(n1060), .CLK(clk_in), .RSTB(n7301), .Q(
        \FIFO[109][17] ) );
  DFFARX1 \FIFO_reg[109][16]  ( .D(n1059), .CLK(clk_in), .RSTB(n7301), .Q(
        \FIFO[109][16] ) );
  DFFARX1 \FIFO_reg[109][15]  ( .D(n1058), .CLK(clk_in), .RSTB(n7301), .Q(
        \FIFO[109][15] ) );
  DFFARX1 \FIFO_reg[109][14]  ( .D(n1057), .CLK(clk_in), .RSTB(n7301), .Q(
        \FIFO[109][14] ) );
  DFFARX1 \FIFO_reg[109][13]  ( .D(n1056), .CLK(clk_in), .RSTB(n7301), .Q(
        \FIFO[109][13] ) );
  DFFARX1 \FIFO_reg[109][12]  ( .D(n1055), .CLK(clk_in), .RSTB(n7301), .Q(
        \FIFO[109][12] ) );
  DFFARX1 \FIFO_reg[109][11]  ( .D(n1054), .CLK(clk_in), .RSTB(n7301), .Q(
        \FIFO[109][11] ) );
  DFFARX1 \FIFO_reg[109][10]  ( .D(n1053), .CLK(clk_in), .RSTB(n7301), .Q(
        \FIFO[109][10] ) );
  DFFARX1 \FIFO_reg[109][9]  ( .D(n1052), .CLK(clk_in), .RSTB(n7301), .Q(
        \FIFO[109][9] ) );
  DFFARX1 \FIFO_reg[109][8]  ( .D(n1051), .CLK(clk_in), .RSTB(n7301), .Q(
        \FIFO[109][8] ) );
  DFFARX1 \FIFO_reg[109][7]  ( .D(n1050), .CLK(clk_in), .RSTB(n7301), .Q(
        \FIFO[109][7] ) );
  DFFARX1 \FIFO_reg[109][6]  ( .D(n1049), .CLK(clk_in), .RSTB(n7301), .Q(
        \FIFO[109][6] ) );
  DFFARX1 \FIFO_reg[109][5]  ( .D(n1048), .CLK(clk_in), .RSTB(n7301), .Q(
        \FIFO[109][5] ) );
  DFFARX1 \FIFO_reg[109][4]  ( .D(n1047), .CLK(clk_in), .RSTB(n7301), .Q(
        \FIFO[109][4] ) );
  DFFARX1 \FIFO_reg[109][3]  ( .D(n1046), .CLK(clk_in), .RSTB(n7302), .Q(
        \FIFO[109][3] ) );
  DFFARX1 \FIFO_reg[109][2]  ( .D(n1045), .CLK(clk_in), .RSTB(n7302), .Q(
        \FIFO[109][2] ) );
  DFFARX1 \FIFO_reg[109][1]  ( .D(n1044), .CLK(clk_in), .RSTB(n7302), .Q(
        \FIFO[109][1] ) );
  DFFARX1 \FIFO_reg[109][0]  ( .D(n1043), .CLK(clk_in), .RSTB(n7302), .Q(
        \FIFO[109][0] ) );
  DFFARX1 \FIFO_reg[110][31]  ( .D(n1042), .CLK(clk_in), .RSTB(n7302), .Q(
        \FIFO[110][31] ) );
  DFFARX1 \FIFO_reg[110][30]  ( .D(n1041), .CLK(clk_in), .RSTB(n7302), .Q(
        \FIFO[110][30] ) );
  DFFARX1 \FIFO_reg[110][29]  ( .D(n1040), .CLK(clk_in), .RSTB(n7302), .Q(
        \FIFO[110][29] ) );
  DFFARX1 \FIFO_reg[110][28]  ( .D(n1039), .CLK(clk_in), .RSTB(n7302), .Q(
        \FIFO[110][28] ) );
  DFFARX1 \FIFO_reg[110][27]  ( .D(n1038), .CLK(clk_in), .RSTB(n7302), .Q(
        \FIFO[110][27] ) );
  DFFARX1 \FIFO_reg[110][26]  ( .D(n1037), .CLK(clk_in), .RSTB(n7302), .Q(
        \FIFO[110][26] ) );
  DFFARX1 \FIFO_reg[110][25]  ( .D(n1036), .CLK(clk_in), .RSTB(n7302), .Q(
        \FIFO[110][25] ) );
  DFFARX1 \FIFO_reg[110][24]  ( .D(n1035), .CLK(clk_in), .RSTB(n7302), .Q(
        \FIFO[110][24] ) );
  DFFARX1 \FIFO_reg[110][23]  ( .D(n1034), .CLK(clk_in), .RSTB(n7302), .Q(
        \FIFO[110][23] ) );
  DFFARX1 \FIFO_reg[110][22]  ( .D(n1033), .CLK(clk_in), .RSTB(n7302), .Q(
        \FIFO[110][22] ) );
  DFFARX1 \FIFO_reg[110][21]  ( .D(n1032), .CLK(clk_in), .RSTB(n7302), .Q(
        \FIFO[110][21] ) );
  DFFARX1 \FIFO_reg[110][20]  ( .D(n1031), .CLK(clk_in), .RSTB(n7302), .Q(
        \FIFO[110][20] ) );
  DFFARX1 \FIFO_reg[110][19]  ( .D(n1030), .CLK(clk_in), .RSTB(n7302), .Q(
        \FIFO[110][19] ) );
  DFFARX1 \FIFO_reg[110][18]  ( .D(n1029), .CLK(clk_in), .RSTB(n7302), .Q(
        \FIFO[110][18] ) );
  DFFARX1 \FIFO_reg[110][17]  ( .D(n1028), .CLK(clk_in), .RSTB(n7303), .Q(
        \FIFO[110][17] ) );
  DFFARX1 \FIFO_reg[110][16]  ( .D(n1027), .CLK(clk_in), .RSTB(n7303), .Q(
        \FIFO[110][16] ) );
  DFFARX1 \FIFO_reg[110][15]  ( .D(n1026), .CLK(clk_in), .RSTB(n7303), .Q(
        \FIFO[110][15] ) );
  DFFARX1 \FIFO_reg[110][14]  ( .D(n1025), .CLK(clk_in), .RSTB(n7303), .Q(
        \FIFO[110][14] ) );
  DFFARX1 \FIFO_reg[110][13]  ( .D(n1024), .CLK(clk_in), .RSTB(n7303), .Q(
        \FIFO[110][13] ) );
  DFFARX1 \FIFO_reg[110][12]  ( .D(n1023), .CLK(clk_in), .RSTB(n7303), .Q(
        \FIFO[110][12] ) );
  DFFARX1 \FIFO_reg[110][11]  ( .D(n1022), .CLK(clk_in), .RSTB(n7303), .Q(
        \FIFO[110][11] ) );
  DFFARX1 \FIFO_reg[110][10]  ( .D(n1021), .CLK(clk_in), .RSTB(n7303), .Q(
        \FIFO[110][10] ) );
  DFFARX1 \FIFO_reg[110][9]  ( .D(n1020), .CLK(clk_in), .RSTB(n7303), .Q(
        \FIFO[110][9] ) );
  DFFARX1 \FIFO_reg[110][8]  ( .D(n1019), .CLK(clk_in), .RSTB(n7303), .Q(
        \FIFO[110][8] ) );
  DFFARX1 \FIFO_reg[110][7]  ( .D(n1018), .CLK(clk_in), .RSTB(n7303), .Q(
        \FIFO[110][7] ) );
  DFFARX1 \FIFO_reg[110][6]  ( .D(n1017), .CLK(clk_in), .RSTB(n7303), .Q(
        \FIFO[110][6] ) );
  DFFARX1 \FIFO_reg[110][5]  ( .D(n1016), .CLK(clk_in), .RSTB(n7303), .Q(
        \FIFO[110][5] ) );
  DFFARX1 \FIFO_reg[110][4]  ( .D(n1015), .CLK(clk_in), .RSTB(n7303), .Q(
        \FIFO[110][4] ) );
  DFFARX1 \FIFO_reg[110][3]  ( .D(n1014), .CLK(clk_in), .RSTB(n7303), .Q(
        \FIFO[110][3] ) );
  DFFARX1 \FIFO_reg[110][2]  ( .D(n1013), .CLK(clk_in), .RSTB(n7303), .Q(
        \FIFO[110][2] ) );
  DFFARX1 \FIFO_reg[110][1]  ( .D(n1012), .CLK(clk_in), .RSTB(n7303), .Q(
        \FIFO[110][1] ) );
  DFFARX1 \FIFO_reg[110][0]  ( .D(n1011), .CLK(clk_in), .RSTB(n7303), .Q(
        \FIFO[110][0] ) );
  DFFARX1 \FIFO_reg[111][31]  ( .D(n1010), .CLK(clk_in), .RSTB(n7304), .Q(
        \FIFO[111][31] ) );
  DFFARX1 \FIFO_reg[111][30]  ( .D(n1009), .CLK(clk_in), .RSTB(n7304), .Q(
        \FIFO[111][30] ) );
  DFFARX1 \FIFO_reg[111][29]  ( .D(n1008), .CLK(clk_in), .RSTB(n7304), .Q(
        \FIFO[111][29] ) );
  DFFARX1 \FIFO_reg[111][28]  ( .D(n1007), .CLK(clk_in), .RSTB(n7304), .Q(
        \FIFO[111][28] ) );
  DFFARX1 \FIFO_reg[111][27]  ( .D(n1006), .CLK(clk_in), .RSTB(n7304), .Q(
        \FIFO[111][27] ) );
  DFFARX1 \FIFO_reg[111][26]  ( .D(n1005), .CLK(clk_in), .RSTB(n7304), .Q(
        \FIFO[111][26] ) );
  DFFARX1 \FIFO_reg[111][25]  ( .D(n1004), .CLK(clk_in), .RSTB(n7304), .Q(
        \FIFO[111][25] ) );
  DFFARX1 \FIFO_reg[111][24]  ( .D(n1003), .CLK(clk_in), .RSTB(n7304), .Q(
        \FIFO[111][24] ) );
  DFFARX1 \FIFO_reg[111][23]  ( .D(n1002), .CLK(clk_in), .RSTB(n7304), .Q(
        \FIFO[111][23] ) );
  DFFARX1 \FIFO_reg[111][22]  ( .D(n1001), .CLK(clk_in), .RSTB(n7304), .Q(
        \FIFO[111][22] ) );
  DFFARX1 \FIFO_reg[111][21]  ( .D(n1000), .CLK(clk_in), .RSTB(n7304), .Q(
        \FIFO[111][21] ) );
  DFFARX1 \FIFO_reg[111][20]  ( .D(n999), .CLK(clk_in), .RSTB(n7304), .Q(
        \FIFO[111][20] ) );
  DFFARX1 \FIFO_reg[111][19]  ( .D(n998), .CLK(clk_in), .RSTB(n7304), .Q(
        \FIFO[111][19] ) );
  DFFARX1 \FIFO_reg[111][18]  ( .D(n997), .CLK(clk_in), .RSTB(n7304), .Q(
        \FIFO[111][18] ) );
  DFFARX1 \FIFO_reg[111][17]  ( .D(n996), .CLK(clk_in), .RSTB(n7304), .Q(
        \FIFO[111][17] ) );
  DFFARX1 \FIFO_reg[111][16]  ( .D(n995), .CLK(clk_in), .RSTB(n7304), .Q(
        \FIFO[111][16] ) );
  DFFARX1 \FIFO_reg[111][15]  ( .D(n994), .CLK(clk_in), .RSTB(n7304), .Q(
        \FIFO[111][15] ) );
  DFFARX1 \FIFO_reg[111][14]  ( .D(n993), .CLK(clk_in), .RSTB(n7304), .Q(
        \FIFO[111][14] ) );
  DFFARX1 \FIFO_reg[111][13]  ( .D(n992), .CLK(clk_in), .RSTB(n7305), .Q(
        \FIFO[111][13] ) );
  DFFARX1 \FIFO_reg[111][12]  ( .D(n991), .CLK(clk_in), .RSTB(n7305), .Q(
        \FIFO[111][12] ) );
  DFFARX1 \FIFO_reg[111][11]  ( .D(n990), .CLK(clk_in), .RSTB(n7305), .Q(
        \FIFO[111][11] ) );
  DFFARX1 \FIFO_reg[111][10]  ( .D(n989), .CLK(clk_in), .RSTB(n7305), .Q(
        \FIFO[111][10] ) );
  DFFARX1 \FIFO_reg[111][9]  ( .D(n988), .CLK(clk_in), .RSTB(n7305), .Q(
        \FIFO[111][9] ) );
  DFFARX1 \FIFO_reg[111][8]  ( .D(n987), .CLK(clk_in), .RSTB(n7305), .Q(
        \FIFO[111][8] ) );
  DFFARX1 \FIFO_reg[111][7]  ( .D(n986), .CLK(clk_in), .RSTB(n7305), .Q(
        \FIFO[111][7] ) );
  DFFARX1 \FIFO_reg[111][6]  ( .D(n985), .CLK(clk_in), .RSTB(n7305), .Q(
        \FIFO[111][6] ) );
  DFFARX1 \FIFO_reg[111][5]  ( .D(n984), .CLK(clk_in), .RSTB(n7305), .Q(
        \FIFO[111][5] ) );
  DFFARX1 \FIFO_reg[111][4]  ( .D(n983), .CLK(clk_in), .RSTB(n7305), .Q(
        \FIFO[111][4] ) );
  DFFARX1 \FIFO_reg[111][3]  ( .D(n982), .CLK(clk_in), .RSTB(n7305), .Q(
        \FIFO[111][3] ) );
  DFFARX1 \FIFO_reg[111][2]  ( .D(n981), .CLK(clk_in), .RSTB(n7305), .Q(
        \FIFO[111][2] ) );
  DFFARX1 \FIFO_reg[111][1]  ( .D(n980), .CLK(clk_in), .RSTB(n7305), .Q(
        \FIFO[111][1] ) );
  DFFARX1 \FIFO_reg[111][0]  ( .D(n979), .CLK(clk_in), .RSTB(n7305), .Q(
        \FIFO[111][0] ) );
  DFFARX1 \FIFO_reg[112][31]  ( .D(n978), .CLK(clk_in), .RSTB(n7305), .Q(
        \FIFO[112][31] ) );
  DFFARX1 \FIFO_reg[112][30]  ( .D(n977), .CLK(clk_in), .RSTB(n7305), .Q(
        \FIFO[112][30] ) );
  DFFARX1 \FIFO_reg[112][29]  ( .D(n976), .CLK(clk_in), .RSTB(n7305), .Q(
        \FIFO[112][29] ) );
  DFFARX1 \FIFO_reg[112][28]  ( .D(n975), .CLK(clk_in), .RSTB(n7305), .Q(
        \FIFO[112][28] ) );
  DFFARX1 \FIFO_reg[112][27]  ( .D(n974), .CLK(clk_in), .RSTB(n7306), .Q(
        \FIFO[112][27] ) );
  DFFARX1 \FIFO_reg[112][26]  ( .D(n973), .CLK(clk_in), .RSTB(n7306), .Q(
        \FIFO[112][26] ) );
  DFFARX1 \FIFO_reg[112][25]  ( .D(n972), .CLK(clk_in), .RSTB(n7306), .Q(
        \FIFO[112][25] ) );
  DFFARX1 \FIFO_reg[112][24]  ( .D(n971), .CLK(clk_in), .RSTB(n7306), .Q(
        \FIFO[112][24] ) );
  DFFARX1 \FIFO_reg[112][23]  ( .D(n970), .CLK(clk_in), .RSTB(n7306), .Q(
        \FIFO[112][23] ) );
  DFFARX1 \FIFO_reg[112][22]  ( .D(n969), .CLK(clk_in), .RSTB(n7306), .Q(
        \FIFO[112][22] ) );
  DFFARX1 \FIFO_reg[112][21]  ( .D(n968), .CLK(clk_in), .RSTB(n7306), .Q(
        \FIFO[112][21] ) );
  DFFARX1 \FIFO_reg[112][20]  ( .D(n967), .CLK(clk_in), .RSTB(n7306), .Q(
        \FIFO[112][20] ) );
  DFFARX1 \FIFO_reg[112][19]  ( .D(n966), .CLK(clk_in), .RSTB(n7306), .Q(
        \FIFO[112][19] ) );
  DFFARX1 \FIFO_reg[112][18]  ( .D(n965), .CLK(clk_in), .RSTB(n7306), .Q(
        \FIFO[112][18] ) );
  DFFARX1 \FIFO_reg[112][17]  ( .D(n964), .CLK(clk_in), .RSTB(n7306), .Q(
        \FIFO[112][17] ) );
  DFFARX1 \FIFO_reg[112][16]  ( .D(n963), .CLK(clk_in), .RSTB(n7306), .Q(
        \FIFO[112][16] ) );
  DFFARX1 \FIFO_reg[112][15]  ( .D(n962), .CLK(clk_in), .RSTB(n7306), .Q(
        \FIFO[112][15] ) );
  DFFARX1 \FIFO_reg[112][14]  ( .D(n961), .CLK(clk_in), .RSTB(n7306), .Q(
        \FIFO[112][14] ) );
  DFFARX1 \FIFO_reg[112][13]  ( .D(n960), .CLK(clk_in), .RSTB(n7306), .Q(
        \FIFO[112][13] ) );
  DFFARX1 \FIFO_reg[112][12]  ( .D(n959), .CLK(clk_in), .RSTB(n7306), .Q(
        \FIFO[112][12] ) );
  DFFARX1 \FIFO_reg[112][11]  ( .D(n958), .CLK(clk_in), .RSTB(n7306), .Q(
        \FIFO[112][11] ) );
  DFFARX1 \FIFO_reg[112][10]  ( .D(n957), .CLK(clk_in), .RSTB(n7306), .Q(
        \FIFO[112][10] ) );
  DFFARX1 \FIFO_reg[112][9]  ( .D(n956), .CLK(clk_in), .RSTB(n7307), .Q(
        \FIFO[112][9] ) );
  DFFARX1 \FIFO_reg[112][8]  ( .D(n955), .CLK(clk_in), .RSTB(n7307), .Q(
        \FIFO[112][8] ) );
  DFFARX1 \FIFO_reg[112][7]  ( .D(n954), .CLK(clk_in), .RSTB(n7307), .Q(
        \FIFO[112][7] ) );
  DFFARX1 \FIFO_reg[112][6]  ( .D(n953), .CLK(clk_in), .RSTB(n7307), .Q(
        \FIFO[112][6] ) );
  DFFARX1 \FIFO_reg[112][5]  ( .D(n952), .CLK(clk_in), .RSTB(n7307), .Q(
        \FIFO[112][5] ) );
  DFFARX1 \FIFO_reg[112][4]  ( .D(n951), .CLK(clk_in), .RSTB(n7307), .Q(
        \FIFO[112][4] ) );
  DFFARX1 \FIFO_reg[112][3]  ( .D(n950), .CLK(clk_in), .RSTB(n7307), .Q(
        \FIFO[112][3] ) );
  DFFARX1 \FIFO_reg[112][2]  ( .D(n949), .CLK(clk_in), .RSTB(n7307), .Q(
        \FIFO[112][2] ) );
  DFFARX1 \FIFO_reg[112][1]  ( .D(n948), .CLK(clk_in), .RSTB(n7307), .Q(
        \FIFO[112][1] ) );
  DFFARX1 \FIFO_reg[112][0]  ( .D(n947), .CLK(clk_in), .RSTB(n7307), .Q(
        \FIFO[112][0] ) );
  DFFARX1 \FIFO_reg[113][31]  ( .D(n946), .CLK(clk_in), .RSTB(n7307), .Q(
        \FIFO[113][31] ) );
  DFFARX1 \FIFO_reg[113][30]  ( .D(n945), .CLK(clk_in), .RSTB(n7307), .Q(
        \FIFO[113][30] ) );
  DFFARX1 \FIFO_reg[113][29]  ( .D(n944), .CLK(clk_in), .RSTB(n7307), .Q(
        \FIFO[113][29] ) );
  DFFARX1 \FIFO_reg[113][28]  ( .D(n943), .CLK(clk_in), .RSTB(n7307), .Q(
        \FIFO[113][28] ) );
  DFFARX1 \FIFO_reg[113][27]  ( .D(n942), .CLK(clk_in), .RSTB(n7307), .Q(
        \FIFO[113][27] ) );
  DFFARX1 \FIFO_reg[113][26]  ( .D(n941), .CLK(clk_in), .RSTB(n7307), .Q(
        \FIFO[113][26] ) );
  DFFARX1 \FIFO_reg[113][25]  ( .D(n940), .CLK(clk_in), .RSTB(n7307), .Q(
        \FIFO[113][25] ) );
  DFFARX1 \FIFO_reg[113][24]  ( .D(n939), .CLK(clk_in), .RSTB(n7307), .Q(
        \FIFO[113][24] ) );
  DFFARX1 \FIFO_reg[113][23]  ( .D(n938), .CLK(clk_in), .RSTB(n7308), .Q(
        \FIFO[113][23] ) );
  DFFARX1 \FIFO_reg[113][22]  ( .D(n937), .CLK(clk_in), .RSTB(n7308), .Q(
        \FIFO[113][22] ) );
  DFFARX1 \FIFO_reg[113][21]  ( .D(n936), .CLK(clk_in), .RSTB(n7308), .Q(
        \FIFO[113][21] ) );
  DFFARX1 \FIFO_reg[113][20]  ( .D(n935), .CLK(clk_in), .RSTB(n7308), .Q(
        \FIFO[113][20] ) );
  DFFARX1 \FIFO_reg[113][19]  ( .D(n934), .CLK(clk_in), .RSTB(n7308), .Q(
        \FIFO[113][19] ) );
  DFFARX1 \FIFO_reg[113][18]  ( .D(n933), .CLK(clk_in), .RSTB(n7308), .Q(
        \FIFO[113][18] ) );
  DFFARX1 \FIFO_reg[113][17]  ( .D(n932), .CLK(clk_in), .RSTB(n7308), .Q(
        \FIFO[113][17] ) );
  DFFARX1 \FIFO_reg[113][16]  ( .D(n931), .CLK(clk_in), .RSTB(n7308), .Q(
        \FIFO[113][16] ) );
  DFFARX1 \FIFO_reg[113][15]  ( .D(n930), .CLK(clk_in), .RSTB(n7308), .Q(
        \FIFO[113][15] ) );
  DFFARX1 \FIFO_reg[113][14]  ( .D(n929), .CLK(clk_in), .RSTB(n7308), .Q(
        \FIFO[113][14] ) );
  DFFARX1 \FIFO_reg[113][13]  ( .D(n928), .CLK(clk_in), .RSTB(n7308), .Q(
        \FIFO[113][13] ) );
  DFFARX1 \FIFO_reg[113][12]  ( .D(n927), .CLK(clk_in), .RSTB(n7308), .Q(
        \FIFO[113][12] ) );
  DFFARX1 \FIFO_reg[113][11]  ( .D(n926), .CLK(clk_in), .RSTB(n7308), .Q(
        \FIFO[113][11] ) );
  DFFARX1 \FIFO_reg[113][10]  ( .D(n925), .CLK(clk_in), .RSTB(n7308), .Q(
        \FIFO[113][10] ) );
  DFFARX1 \FIFO_reg[113][9]  ( .D(n924), .CLK(clk_in), .RSTB(n7308), .Q(
        \FIFO[113][9] ) );
  DFFARX1 \FIFO_reg[113][8]  ( .D(n923), .CLK(clk_in), .RSTB(n7308), .Q(
        \FIFO[113][8] ) );
  DFFARX1 \FIFO_reg[113][7]  ( .D(n922), .CLK(clk_in), .RSTB(n7308), .Q(
        \FIFO[113][7] ) );
  DFFARX1 \FIFO_reg[113][6]  ( .D(n921), .CLK(clk_in), .RSTB(n7308), .Q(
        \FIFO[113][6] ) );
  DFFARX1 \FIFO_reg[113][5]  ( .D(n920), .CLK(clk_in), .RSTB(n7309), .Q(
        \FIFO[113][5] ) );
  DFFARX1 \FIFO_reg[113][4]  ( .D(n919), .CLK(clk_in), .RSTB(n7309), .Q(
        \FIFO[113][4] ) );
  DFFARX1 \FIFO_reg[113][3]  ( .D(n918), .CLK(clk_in), .RSTB(n7309), .Q(
        \FIFO[113][3] ) );
  DFFARX1 \FIFO_reg[113][2]  ( .D(n917), .CLK(clk_in), .RSTB(n7309), .Q(
        \FIFO[113][2] ) );
  DFFARX1 \FIFO_reg[113][1]  ( .D(n916), .CLK(clk_in), .RSTB(n7309), .Q(
        \FIFO[113][1] ) );
  DFFARX1 \FIFO_reg[113][0]  ( .D(n915), .CLK(clk_in), .RSTB(n7309), .Q(
        \FIFO[113][0] ) );
  DFFARX1 \FIFO_reg[114][31]  ( .D(n914), .CLK(clk_in), .RSTB(n7309), .Q(
        \FIFO[114][31] ) );
  DFFARX1 \FIFO_reg[114][30]  ( .D(n913), .CLK(clk_in), .RSTB(n7309), .Q(
        \FIFO[114][30] ) );
  DFFARX1 \FIFO_reg[114][29]  ( .D(n912), .CLK(clk_in), .RSTB(n7309), .Q(
        \FIFO[114][29] ) );
  DFFARX1 \FIFO_reg[114][28]  ( .D(n911), .CLK(clk_in), .RSTB(n7309), .Q(
        \FIFO[114][28] ) );
  DFFARX1 \FIFO_reg[114][27]  ( .D(n910), .CLK(clk_in), .RSTB(n7309), .Q(
        \FIFO[114][27] ) );
  DFFARX1 \FIFO_reg[114][26]  ( .D(n909), .CLK(clk_in), .RSTB(n7309), .Q(
        \FIFO[114][26] ) );
  DFFARX1 \FIFO_reg[114][25]  ( .D(n908), .CLK(clk_in), .RSTB(n7309), .Q(
        \FIFO[114][25] ) );
  DFFARX1 \FIFO_reg[114][24]  ( .D(n907), .CLK(clk_in), .RSTB(n7309), .Q(
        \FIFO[114][24] ) );
  DFFARX1 \FIFO_reg[114][23]  ( .D(n906), .CLK(clk_in), .RSTB(n7309), .Q(
        \FIFO[114][23] ) );
  DFFARX1 \FIFO_reg[114][22]  ( .D(n905), .CLK(clk_in), .RSTB(n7309), .Q(
        \FIFO[114][22] ) );
  DFFARX1 \FIFO_reg[114][21]  ( .D(n904), .CLK(clk_in), .RSTB(n7309), .Q(
        \FIFO[114][21] ) );
  DFFARX1 \FIFO_reg[114][20]  ( .D(n903), .CLK(clk_in), .RSTB(n7309), .Q(
        \FIFO[114][20] ) );
  DFFARX1 \FIFO_reg[114][19]  ( .D(n902), .CLK(clk_in), .RSTB(n7310), .Q(
        \FIFO[114][19] ) );
  DFFARX1 \FIFO_reg[114][18]  ( .D(n901), .CLK(clk_in), .RSTB(n7310), .Q(
        \FIFO[114][18] ) );
  DFFARX1 \FIFO_reg[114][17]  ( .D(n900), .CLK(clk_in), .RSTB(n7310), .Q(
        \FIFO[114][17] ) );
  DFFARX1 \FIFO_reg[114][16]  ( .D(n899), .CLK(clk_in), .RSTB(n7310), .Q(
        \FIFO[114][16] ) );
  DFFARX1 \FIFO_reg[114][15]  ( .D(n898), .CLK(clk_in), .RSTB(n7310), .Q(
        \FIFO[114][15] ) );
  DFFARX1 \FIFO_reg[114][14]  ( .D(n897), .CLK(clk_in), .RSTB(n7310), .Q(
        \FIFO[114][14] ) );
  DFFARX1 \FIFO_reg[114][13]  ( .D(n896), .CLK(clk_in), .RSTB(n7310), .Q(
        \FIFO[114][13] ) );
  DFFARX1 \FIFO_reg[114][12]  ( .D(n895), .CLK(clk_in), .RSTB(n7310), .Q(
        \FIFO[114][12] ) );
  DFFARX1 \FIFO_reg[114][11]  ( .D(n894), .CLK(clk_in), .RSTB(n7310), .Q(
        \FIFO[114][11] ) );
  DFFARX1 \FIFO_reg[114][10]  ( .D(n893), .CLK(clk_in), .RSTB(n7310), .Q(
        \FIFO[114][10] ) );
  DFFARX1 \FIFO_reg[114][9]  ( .D(n892), .CLK(clk_in), .RSTB(n7310), .Q(
        \FIFO[114][9] ) );
  DFFARX1 \FIFO_reg[114][8]  ( .D(n891), .CLK(clk_in), .RSTB(n7310), .Q(
        \FIFO[114][8] ) );
  DFFARX1 \FIFO_reg[114][7]  ( .D(n890), .CLK(clk_in), .RSTB(n7310), .Q(
        \FIFO[114][7] ) );
  DFFARX1 \FIFO_reg[114][6]  ( .D(n889), .CLK(clk_in), .RSTB(n7310), .Q(
        \FIFO[114][6] ) );
  DFFARX1 \FIFO_reg[114][5]  ( .D(n888), .CLK(clk_in), .RSTB(n7310), .Q(
        \FIFO[114][5] ) );
  DFFARX1 \FIFO_reg[114][4]  ( .D(n887), .CLK(clk_in), .RSTB(n7310), .Q(
        \FIFO[114][4] ) );
  DFFARX1 \FIFO_reg[114][3]  ( .D(n886), .CLK(clk_in), .RSTB(n7310), .Q(
        \FIFO[114][3] ) );
  DFFARX1 \FIFO_reg[114][2]  ( .D(n885), .CLK(clk_in), .RSTB(n7310), .Q(
        \FIFO[114][2] ) );
  DFFARX1 \FIFO_reg[114][1]  ( .D(n884), .CLK(clk_in), .RSTB(n7311), .Q(
        \FIFO[114][1] ) );
  DFFARX1 \FIFO_reg[114][0]  ( .D(n883), .CLK(clk_in), .RSTB(n7311), .Q(
        \FIFO[114][0] ) );
  DFFARX1 \FIFO_reg[115][31]  ( .D(n882), .CLK(clk_in), .RSTB(n7311), .Q(
        \FIFO[115][31] ) );
  DFFARX1 \FIFO_reg[115][30]  ( .D(n881), .CLK(clk_in), .RSTB(n7311), .Q(
        \FIFO[115][30] ) );
  DFFARX1 \FIFO_reg[115][29]  ( .D(n880), .CLK(clk_in), .RSTB(n7311), .Q(
        \FIFO[115][29] ) );
  DFFARX1 \FIFO_reg[115][28]  ( .D(n879), .CLK(clk_in), .RSTB(n7311), .Q(
        \FIFO[115][28] ) );
  DFFARX1 \FIFO_reg[115][27]  ( .D(n878), .CLK(clk_in), .RSTB(n7311), .Q(
        \FIFO[115][27] ) );
  DFFARX1 \FIFO_reg[115][26]  ( .D(n877), .CLK(clk_in), .RSTB(n7311), .Q(
        \FIFO[115][26] ) );
  DFFARX1 \FIFO_reg[115][25]  ( .D(n876), .CLK(clk_in), .RSTB(n7311), .Q(
        \FIFO[115][25] ) );
  DFFARX1 \FIFO_reg[115][24]  ( .D(n875), .CLK(clk_in), .RSTB(n7311), .Q(
        \FIFO[115][24] ) );
  DFFARX1 \FIFO_reg[115][23]  ( .D(n874), .CLK(clk_in), .RSTB(n7311), .Q(
        \FIFO[115][23] ) );
  DFFARX1 \FIFO_reg[115][22]  ( .D(n873), .CLK(clk_in), .RSTB(n7311), .Q(
        \FIFO[115][22] ) );
  DFFARX1 \FIFO_reg[115][21]  ( .D(n872), .CLK(clk_in), .RSTB(n7311), .Q(
        \FIFO[115][21] ) );
  DFFARX1 \FIFO_reg[115][20]  ( .D(n871), .CLK(clk_in), .RSTB(n7311), .Q(
        \FIFO[115][20] ) );
  DFFARX1 \FIFO_reg[115][19]  ( .D(n870), .CLK(clk_in), .RSTB(n7311), .Q(
        \FIFO[115][19] ) );
  DFFARX1 \FIFO_reg[115][18]  ( .D(n869), .CLK(clk_in), .RSTB(n7311), .Q(
        \FIFO[115][18] ) );
  DFFARX1 \FIFO_reg[115][17]  ( .D(n868), .CLK(clk_in), .RSTB(n7311), .Q(
        \FIFO[115][17] ) );
  DFFARX1 \FIFO_reg[115][16]  ( .D(n867), .CLK(clk_in), .RSTB(n7311), .Q(
        \FIFO[115][16] ) );
  DFFARX1 \FIFO_reg[115][15]  ( .D(n866), .CLK(clk_in), .RSTB(n7312), .Q(
        \FIFO[115][15] ) );
  DFFARX1 \FIFO_reg[115][14]  ( .D(n865), .CLK(clk_in), .RSTB(n7312), .Q(
        \FIFO[115][14] ) );
  DFFARX1 \FIFO_reg[115][13]  ( .D(n864), .CLK(clk_in), .RSTB(n7312), .Q(
        \FIFO[115][13] ) );
  DFFARX1 \FIFO_reg[115][12]  ( .D(n863), .CLK(clk_in), .RSTB(n7312), .Q(
        \FIFO[115][12] ) );
  DFFARX1 \FIFO_reg[115][11]  ( .D(n862), .CLK(clk_in), .RSTB(n7312), .Q(
        \FIFO[115][11] ) );
  DFFARX1 \FIFO_reg[115][10]  ( .D(n861), .CLK(clk_in), .RSTB(n7312), .Q(
        \FIFO[115][10] ) );
  DFFARX1 \FIFO_reg[115][9]  ( .D(n860), .CLK(clk_in), .RSTB(n7312), .Q(
        \FIFO[115][9] ) );
  DFFARX1 \FIFO_reg[115][8]  ( .D(n859), .CLK(clk_in), .RSTB(n7312), .Q(
        \FIFO[115][8] ) );
  DFFARX1 \FIFO_reg[115][7]  ( .D(n858), .CLK(clk_in), .RSTB(n7312), .Q(
        \FIFO[115][7] ) );
  DFFARX1 \FIFO_reg[115][6]  ( .D(n857), .CLK(clk_in), .RSTB(n7312), .Q(
        \FIFO[115][6] ) );
  DFFARX1 \FIFO_reg[115][5]  ( .D(n856), .CLK(clk_in), .RSTB(n7312), .Q(
        \FIFO[115][5] ) );
  DFFARX1 \FIFO_reg[115][4]  ( .D(n855), .CLK(clk_in), .RSTB(n7312), .Q(
        \FIFO[115][4] ) );
  DFFARX1 \FIFO_reg[115][3]  ( .D(n854), .CLK(clk_in), .RSTB(n7312), .Q(
        \FIFO[115][3] ) );
  DFFARX1 \FIFO_reg[115][2]  ( .D(n853), .CLK(clk_in), .RSTB(n7312), .Q(
        \FIFO[115][2] ) );
  DFFARX1 \FIFO_reg[115][1]  ( .D(n852), .CLK(clk_in), .RSTB(n7312), .Q(
        \FIFO[115][1] ) );
  DFFARX1 \FIFO_reg[115][0]  ( .D(n851), .CLK(clk_in), .RSTB(n7312), .Q(
        \FIFO[115][0] ) );
  DFFARX1 \FIFO_reg[116][31]  ( .D(n850), .CLK(clk_in), .RSTB(n7312), .Q(
        \FIFO[116][31] ) );
  DFFARX1 \FIFO_reg[116][30]  ( .D(n849), .CLK(clk_in), .RSTB(n7312), .Q(
        \FIFO[116][30] ) );
  DFFARX1 \FIFO_reg[116][29]  ( .D(n848), .CLK(clk_in), .RSTB(n7313), .Q(
        \FIFO[116][29] ) );
  DFFARX1 \FIFO_reg[116][28]  ( .D(n847), .CLK(clk_in), .RSTB(n7313), .Q(
        \FIFO[116][28] ) );
  DFFARX1 \FIFO_reg[116][27]  ( .D(n846), .CLK(clk_in), .RSTB(n7313), .Q(
        \FIFO[116][27] ) );
  DFFARX1 \FIFO_reg[116][26]  ( .D(n845), .CLK(clk_in), .RSTB(n7313), .Q(
        \FIFO[116][26] ) );
  DFFARX1 \FIFO_reg[116][25]  ( .D(n844), .CLK(clk_in), .RSTB(n7313), .Q(
        \FIFO[116][25] ) );
  DFFARX1 \FIFO_reg[116][24]  ( .D(n843), .CLK(clk_in), .RSTB(n7313), .Q(
        \FIFO[116][24] ) );
  DFFARX1 \FIFO_reg[116][23]  ( .D(n842), .CLK(clk_in), .RSTB(n7313), .Q(
        \FIFO[116][23] ) );
  DFFARX1 \FIFO_reg[116][22]  ( .D(n841), .CLK(clk_in), .RSTB(n7313), .Q(
        \FIFO[116][22] ) );
  DFFARX1 \FIFO_reg[116][21]  ( .D(n840), .CLK(clk_in), .RSTB(n7313), .Q(
        \FIFO[116][21] ) );
  DFFARX1 \FIFO_reg[116][20]  ( .D(n839), .CLK(clk_in), .RSTB(n7313), .Q(
        \FIFO[116][20] ) );
  DFFARX1 \FIFO_reg[116][19]  ( .D(n838), .CLK(clk_in), .RSTB(n7313), .Q(
        \FIFO[116][19] ) );
  DFFARX1 \FIFO_reg[116][18]  ( .D(n837), .CLK(clk_in), .RSTB(n7313), .Q(
        \FIFO[116][18] ) );
  DFFARX1 \FIFO_reg[116][17]  ( .D(n836), .CLK(clk_in), .RSTB(n7313), .Q(
        \FIFO[116][17] ) );
  DFFARX1 \FIFO_reg[116][16]  ( .D(n835), .CLK(clk_in), .RSTB(n7313), .Q(
        \FIFO[116][16] ) );
  DFFARX1 \FIFO_reg[116][15]  ( .D(n834), .CLK(clk_in), .RSTB(n7313), .Q(
        \FIFO[116][15] ) );
  DFFARX1 \FIFO_reg[116][14]  ( .D(n833), .CLK(clk_in), .RSTB(n7313), .Q(
        \FIFO[116][14] ) );
  DFFARX1 \FIFO_reg[116][13]  ( .D(n832), .CLK(clk_in), .RSTB(n7313), .Q(
        \FIFO[116][13] ) );
  DFFARX1 \FIFO_reg[116][12]  ( .D(n831), .CLK(clk_in), .RSTB(n7313), .Q(
        \FIFO[116][12] ) );
  DFFARX1 \FIFO_reg[116][11]  ( .D(n830), .CLK(clk_in), .RSTB(n7314), .Q(
        \FIFO[116][11] ) );
  DFFARX1 \FIFO_reg[116][10]  ( .D(n829), .CLK(clk_in), .RSTB(n7314), .Q(
        \FIFO[116][10] ) );
  DFFARX1 \FIFO_reg[116][9]  ( .D(n828), .CLK(clk_in), .RSTB(n7314), .Q(
        \FIFO[116][9] ) );
  DFFARX1 \FIFO_reg[116][8]  ( .D(n827), .CLK(clk_in), .RSTB(n7314), .Q(
        \FIFO[116][8] ) );
  DFFARX1 \FIFO_reg[116][7]  ( .D(n826), .CLK(clk_in), .RSTB(n7314), .Q(
        \FIFO[116][7] ) );
  DFFARX1 \FIFO_reg[116][6]  ( .D(n825), .CLK(clk_in), .RSTB(n7314), .Q(
        \FIFO[116][6] ) );
  DFFARX1 \FIFO_reg[116][5]  ( .D(n824), .CLK(clk_in), .RSTB(n7314), .Q(
        \FIFO[116][5] ) );
  DFFARX1 \FIFO_reg[116][4]  ( .D(n823), .CLK(clk_in), .RSTB(n7314), .Q(
        \FIFO[116][4] ) );
  DFFARX1 \FIFO_reg[116][3]  ( .D(n822), .CLK(clk_in), .RSTB(n7314), .Q(
        \FIFO[116][3] ) );
  DFFARX1 \FIFO_reg[116][2]  ( .D(n821), .CLK(clk_in), .RSTB(n7314), .Q(
        \FIFO[116][2] ) );
  DFFARX1 \FIFO_reg[116][1]  ( .D(n820), .CLK(clk_in), .RSTB(n7314), .Q(
        \FIFO[116][1] ) );
  DFFARX1 \FIFO_reg[116][0]  ( .D(n819), .CLK(clk_in), .RSTB(n7314), .Q(
        \FIFO[116][0] ) );
  DFFARX1 \FIFO_reg[117][31]  ( .D(n818), .CLK(clk_in), .RSTB(n7314), .Q(
        \FIFO[117][31] ) );
  DFFARX1 \FIFO_reg[117][30]  ( .D(n817), .CLK(clk_in), .RSTB(n7314), .Q(
        \FIFO[117][30] ) );
  DFFARX1 \FIFO_reg[117][29]  ( .D(n816), .CLK(clk_in), .RSTB(n7314), .Q(
        \FIFO[117][29] ) );
  DFFARX1 \FIFO_reg[117][28]  ( .D(n815), .CLK(clk_in), .RSTB(n7314), .Q(
        \FIFO[117][28] ) );
  DFFARX1 \FIFO_reg[117][27]  ( .D(n814), .CLK(clk_in), .RSTB(n7314), .Q(
        \FIFO[117][27] ) );
  DFFARX1 \FIFO_reg[117][26]  ( .D(n813), .CLK(clk_in), .RSTB(n7314), .Q(
        \FIFO[117][26] ) );
  DFFARX1 \FIFO_reg[117][25]  ( .D(n812), .CLK(clk_in), .RSTB(n7315), .Q(
        \FIFO[117][25] ) );
  DFFARX1 \FIFO_reg[117][24]  ( .D(n811), .CLK(clk_in), .RSTB(n7315), .Q(
        \FIFO[117][24] ) );
  DFFARX1 \FIFO_reg[117][23]  ( .D(n810), .CLK(clk_in), .RSTB(n7315), .Q(
        \FIFO[117][23] ) );
  DFFARX1 \FIFO_reg[117][22]  ( .D(n809), .CLK(clk_in), .RSTB(n7315), .Q(
        \FIFO[117][22] ) );
  DFFARX1 \FIFO_reg[117][21]  ( .D(n808), .CLK(clk_in), .RSTB(n7315), .Q(
        \FIFO[117][21] ) );
  DFFARX1 \FIFO_reg[117][20]  ( .D(n807), .CLK(clk_in), .RSTB(n7315), .Q(
        \FIFO[117][20] ) );
  DFFARX1 \FIFO_reg[117][19]  ( .D(n806), .CLK(clk_in), .RSTB(n7315), .Q(
        \FIFO[117][19] ) );
  DFFARX1 \FIFO_reg[117][18]  ( .D(n805), .CLK(clk_in), .RSTB(n7315), .Q(
        \FIFO[117][18] ) );
  DFFARX1 \FIFO_reg[117][17]  ( .D(n804), .CLK(clk_in), .RSTB(n7315), .Q(
        \FIFO[117][17] ) );
  DFFARX1 \FIFO_reg[117][16]  ( .D(n803), .CLK(clk_in), .RSTB(n7315), .Q(
        \FIFO[117][16] ) );
  DFFARX1 \FIFO_reg[117][15]  ( .D(n802), .CLK(clk_in), .RSTB(n7315), .Q(
        \FIFO[117][15] ) );
  DFFARX1 \FIFO_reg[117][14]  ( .D(n801), .CLK(clk_in), .RSTB(n7315), .Q(
        \FIFO[117][14] ) );
  DFFARX1 \FIFO_reg[117][13]  ( .D(n800), .CLK(clk_in), .RSTB(n7315), .Q(
        \FIFO[117][13] ) );
  DFFARX1 \FIFO_reg[117][12]  ( .D(n799), .CLK(clk_in), .RSTB(n7315), .Q(
        \FIFO[117][12] ) );
  DFFARX1 \FIFO_reg[117][11]  ( .D(n798), .CLK(clk_in), .RSTB(n7315), .Q(
        \FIFO[117][11] ) );
  DFFARX1 \FIFO_reg[117][10]  ( .D(n797), .CLK(clk_in), .RSTB(n7315), .Q(
        \FIFO[117][10] ) );
  DFFARX1 \FIFO_reg[117][9]  ( .D(n796), .CLK(clk_in), .RSTB(n7315), .Q(
        \FIFO[117][9] ) );
  DFFARX1 \FIFO_reg[117][8]  ( .D(n795), .CLK(clk_in), .RSTB(n7315), .Q(
        \FIFO[117][8] ) );
  DFFARX1 \FIFO_reg[117][7]  ( .D(n794), .CLK(clk_in), .RSTB(n7316), .Q(
        \FIFO[117][7] ) );
  DFFARX1 \FIFO_reg[117][6]  ( .D(n793), .CLK(clk_in), .RSTB(n7316), .Q(
        \FIFO[117][6] ) );
  DFFARX1 \FIFO_reg[117][5]  ( .D(n792), .CLK(clk_in), .RSTB(n7316), .Q(
        \FIFO[117][5] ) );
  DFFARX1 \FIFO_reg[117][4]  ( .D(n791), .CLK(clk_in), .RSTB(n7316), .Q(
        \FIFO[117][4] ) );
  DFFARX1 \FIFO_reg[117][3]  ( .D(n790), .CLK(clk_in), .RSTB(n7316), .Q(
        \FIFO[117][3] ) );
  DFFARX1 \FIFO_reg[117][2]  ( .D(n789), .CLK(clk_in), .RSTB(n7316), .Q(
        \FIFO[117][2] ) );
  DFFARX1 \FIFO_reg[117][1]  ( .D(n788), .CLK(clk_in), .RSTB(n7316), .Q(
        \FIFO[117][1] ) );
  DFFARX1 \FIFO_reg[117][0]  ( .D(n787), .CLK(clk_in), .RSTB(n7316), .Q(
        \FIFO[117][0] ) );
  DFFARX1 \FIFO_reg[118][31]  ( .D(n786), .CLK(clk_in), .RSTB(n7316), .Q(
        \FIFO[118][31] ) );
  DFFARX1 \FIFO_reg[118][30]  ( .D(n785), .CLK(clk_in), .RSTB(n7316), .Q(
        \FIFO[118][30] ) );
  DFFARX1 \FIFO_reg[118][29]  ( .D(n784), .CLK(clk_in), .RSTB(n7316), .Q(
        \FIFO[118][29] ) );
  DFFARX1 \FIFO_reg[118][28]  ( .D(n783), .CLK(clk_in), .RSTB(n7316), .Q(
        \FIFO[118][28] ) );
  DFFARX1 \FIFO_reg[118][27]  ( .D(n782), .CLK(clk_in), .RSTB(n7316), .Q(
        \FIFO[118][27] ) );
  DFFARX1 \FIFO_reg[118][26]  ( .D(n781), .CLK(clk_in), .RSTB(n7316), .Q(
        \FIFO[118][26] ) );
  DFFARX1 \FIFO_reg[118][25]  ( .D(n780), .CLK(clk_in), .RSTB(n7316), .Q(
        \FIFO[118][25] ) );
  DFFARX1 \FIFO_reg[118][24]  ( .D(n779), .CLK(clk_in), .RSTB(n7316), .Q(
        \FIFO[118][24] ) );
  DFFARX1 \FIFO_reg[118][23]  ( .D(n778), .CLK(clk_in), .RSTB(n7316), .Q(
        \FIFO[118][23] ) );
  DFFARX1 \FIFO_reg[118][22]  ( .D(n777), .CLK(clk_in), .RSTB(n7316), .Q(
        \FIFO[118][22] ) );
  DFFARX1 \FIFO_reg[118][21]  ( .D(n776), .CLK(clk_in), .RSTB(n7317), .Q(
        \FIFO[118][21] ) );
  DFFARX1 \FIFO_reg[118][20]  ( .D(n775), .CLK(clk_in), .RSTB(n7317), .Q(
        \FIFO[118][20] ) );
  DFFARX1 \FIFO_reg[118][19]  ( .D(n774), .CLK(clk_in), .RSTB(n7317), .Q(
        \FIFO[118][19] ) );
  DFFARX1 \FIFO_reg[118][18]  ( .D(n773), .CLK(clk_in), .RSTB(n7317), .Q(
        \FIFO[118][18] ) );
  DFFARX1 \FIFO_reg[118][17]  ( .D(n772), .CLK(clk_in), .RSTB(n7317), .Q(
        \FIFO[118][17] ) );
  DFFARX1 \FIFO_reg[118][16]  ( .D(n771), .CLK(clk_in), .RSTB(n7317), .Q(
        \FIFO[118][16] ) );
  DFFARX1 \FIFO_reg[118][15]  ( .D(n770), .CLK(clk_in), .RSTB(n7317), .Q(
        \FIFO[118][15] ) );
  DFFARX1 \FIFO_reg[118][14]  ( .D(n769), .CLK(clk_in), .RSTB(n7317), .Q(
        \FIFO[118][14] ) );
  DFFARX1 \FIFO_reg[118][13]  ( .D(n768), .CLK(clk_in), .RSTB(n7317), .Q(
        \FIFO[118][13] ) );
  DFFARX1 \FIFO_reg[118][12]  ( .D(n767), .CLK(clk_in), .RSTB(n7317), .Q(
        \FIFO[118][12] ) );
  DFFARX1 \FIFO_reg[118][11]  ( .D(n766), .CLK(clk_in), .RSTB(n7317), .Q(
        \FIFO[118][11] ) );
  DFFARX1 \FIFO_reg[118][10]  ( .D(n765), .CLK(clk_in), .RSTB(n7317), .Q(
        \FIFO[118][10] ) );
  DFFARX1 \FIFO_reg[118][9]  ( .D(n764), .CLK(clk_in), .RSTB(n7317), .Q(
        \FIFO[118][9] ) );
  DFFARX1 \FIFO_reg[118][8]  ( .D(n763), .CLK(clk_in), .RSTB(n7317), .Q(
        \FIFO[118][8] ) );
  DFFARX1 \FIFO_reg[118][7]  ( .D(n762), .CLK(clk_in), .RSTB(n7317), .Q(
        \FIFO[118][7] ) );
  DFFARX1 \FIFO_reg[118][6]  ( .D(n761), .CLK(clk_in), .RSTB(n7317), .Q(
        \FIFO[118][6] ) );
  DFFARX1 \FIFO_reg[118][5]  ( .D(n760), .CLK(clk_in), .RSTB(n7317), .Q(
        \FIFO[118][5] ) );
  DFFARX1 \FIFO_reg[118][4]  ( .D(n759), .CLK(clk_in), .RSTB(n7317), .Q(
        \FIFO[118][4] ) );
  DFFARX1 \FIFO_reg[118][3]  ( .D(n758), .CLK(clk_in), .RSTB(n7318), .Q(
        \FIFO[118][3] ) );
  DFFARX1 \FIFO_reg[118][2]  ( .D(n757), .CLK(clk_in), .RSTB(n7318), .Q(
        \FIFO[118][2] ) );
  DFFARX1 \FIFO_reg[118][1]  ( .D(n756), .CLK(clk_in), .RSTB(n7318), .Q(
        \FIFO[118][1] ) );
  DFFARX1 \FIFO_reg[118][0]  ( .D(n755), .CLK(clk_in), .RSTB(n7318), .Q(
        \FIFO[118][0] ) );
  DFFARX1 \FIFO_reg[119][31]  ( .D(n754), .CLK(clk_in), .RSTB(n7318), .Q(
        \FIFO[119][31] ) );
  DFFARX1 \FIFO_reg[119][30]  ( .D(n753), .CLK(clk_in), .RSTB(n7318), .Q(
        \FIFO[119][30] ) );
  DFFARX1 \FIFO_reg[119][29]  ( .D(n752), .CLK(clk_in), .RSTB(n7318), .Q(
        \FIFO[119][29] ) );
  DFFARX1 \FIFO_reg[119][28]  ( .D(n751), .CLK(clk_in), .RSTB(n7318), .Q(
        \FIFO[119][28] ) );
  DFFARX1 \FIFO_reg[119][27]  ( .D(n750), .CLK(clk_in), .RSTB(n7318), .Q(
        \FIFO[119][27] ) );
  DFFARX1 \FIFO_reg[119][26]  ( .D(n749), .CLK(clk_in), .RSTB(n7318), .Q(
        \FIFO[119][26] ) );
  DFFARX1 \FIFO_reg[119][25]  ( .D(n748), .CLK(clk_in), .RSTB(n7318), .Q(
        \FIFO[119][25] ) );
  DFFARX1 \FIFO_reg[119][24]  ( .D(n747), .CLK(clk_in), .RSTB(n7318), .Q(
        \FIFO[119][24] ) );
  DFFARX1 \FIFO_reg[119][23]  ( .D(n746), .CLK(clk_in), .RSTB(n7318), .Q(
        \FIFO[119][23] ) );
  DFFARX1 \FIFO_reg[119][22]  ( .D(n745), .CLK(clk_in), .RSTB(n7318), .Q(
        \FIFO[119][22] ) );
  DFFARX1 \FIFO_reg[119][21]  ( .D(n744), .CLK(clk_in), .RSTB(n7318), .Q(
        \FIFO[119][21] ) );
  DFFARX1 \FIFO_reg[119][20]  ( .D(n743), .CLK(clk_in), .RSTB(n7318), .Q(
        \FIFO[119][20] ) );
  DFFARX1 \FIFO_reg[119][19]  ( .D(n742), .CLK(clk_in), .RSTB(n7318), .Q(
        \FIFO[119][19] ) );
  DFFARX1 \FIFO_reg[119][18]  ( .D(n741), .CLK(clk_in), .RSTB(n7318), .Q(
        \FIFO[119][18] ) );
  DFFARX1 \FIFO_reg[119][17]  ( .D(n740), .CLK(clk_in), .RSTB(n7319), .Q(
        \FIFO[119][17] ) );
  DFFARX1 \FIFO_reg[119][16]  ( .D(n739), .CLK(clk_in), .RSTB(n7319), .Q(
        \FIFO[119][16] ) );
  DFFARX1 \FIFO_reg[119][15]  ( .D(n738), .CLK(clk_in), .RSTB(n7319), .Q(
        \FIFO[119][15] ) );
  DFFARX1 \FIFO_reg[119][14]  ( .D(n737), .CLK(clk_in), .RSTB(n7319), .Q(
        \FIFO[119][14] ) );
  DFFARX1 \FIFO_reg[119][13]  ( .D(n736), .CLK(clk_in), .RSTB(n7319), .Q(
        \FIFO[119][13] ) );
  DFFARX1 \FIFO_reg[119][12]  ( .D(n735), .CLK(clk_in), .RSTB(n7319), .Q(
        \FIFO[119][12] ) );
  DFFARX1 \FIFO_reg[119][11]  ( .D(n734), .CLK(clk_in), .RSTB(n7319), .Q(
        \FIFO[119][11] ) );
  DFFARX1 \FIFO_reg[119][10]  ( .D(n733), .CLK(clk_in), .RSTB(n7319), .Q(
        \FIFO[119][10] ) );
  DFFARX1 \FIFO_reg[119][9]  ( .D(n732), .CLK(clk_in), .RSTB(n7319), .Q(
        \FIFO[119][9] ) );
  DFFARX1 \FIFO_reg[119][8]  ( .D(n731), .CLK(clk_in), .RSTB(n7319), .Q(
        \FIFO[119][8] ) );
  DFFARX1 \FIFO_reg[119][7]  ( .D(n730), .CLK(clk_in), .RSTB(n7319), .Q(
        \FIFO[119][7] ) );
  DFFARX1 \FIFO_reg[119][6]  ( .D(n729), .CLK(clk_in), .RSTB(n7319), .Q(
        \FIFO[119][6] ) );
  DFFARX1 \FIFO_reg[119][5]  ( .D(n728), .CLK(clk_in), .RSTB(n7319), .Q(
        \FIFO[119][5] ) );
  DFFARX1 \FIFO_reg[119][4]  ( .D(n727), .CLK(clk_in), .RSTB(n7319), .Q(
        \FIFO[119][4] ) );
  DFFARX1 \FIFO_reg[119][3]  ( .D(n726), .CLK(clk_in), .RSTB(n7319), .Q(
        \FIFO[119][3] ) );
  DFFARX1 \FIFO_reg[119][2]  ( .D(n725), .CLK(clk_in), .RSTB(n7319), .Q(
        \FIFO[119][2] ) );
  DFFARX1 \FIFO_reg[119][1]  ( .D(n724), .CLK(clk_in), .RSTB(n7319), .Q(
        \FIFO[119][1] ) );
  DFFARX1 \FIFO_reg[119][0]  ( .D(n723), .CLK(clk_in), .RSTB(n7319), .Q(
        \FIFO[119][0] ) );
  DFFARX1 \FIFO_reg[120][31]  ( .D(n722), .CLK(clk_in), .RSTB(n7320), .Q(
        \FIFO[120][31] ) );
  DFFARX1 \FIFO_reg[120][30]  ( .D(n721), .CLK(clk_in), .RSTB(n7320), .Q(
        \FIFO[120][30] ) );
  DFFARX1 \FIFO_reg[120][29]  ( .D(n720), .CLK(clk_in), .RSTB(n7320), .Q(
        \FIFO[120][29] ) );
  DFFARX1 \FIFO_reg[120][28]  ( .D(n719), .CLK(clk_in), .RSTB(n7320), .Q(
        \FIFO[120][28] ) );
  DFFARX1 \FIFO_reg[120][27]  ( .D(n718), .CLK(clk_in), .RSTB(n7320), .Q(
        \FIFO[120][27] ) );
  DFFARX1 \FIFO_reg[120][26]  ( .D(n717), .CLK(clk_in), .RSTB(n7320), .Q(
        \FIFO[120][26] ) );
  DFFARX1 \FIFO_reg[120][25]  ( .D(n716), .CLK(clk_in), .RSTB(n7320), .Q(
        \FIFO[120][25] ) );
  DFFARX1 \FIFO_reg[120][24]  ( .D(n715), .CLK(clk_in), .RSTB(n7320), .Q(
        \FIFO[120][24] ) );
  DFFARX1 \FIFO_reg[120][23]  ( .D(n714), .CLK(clk_in), .RSTB(n7320), .Q(
        \FIFO[120][23] ) );
  DFFARX1 \FIFO_reg[120][22]  ( .D(n713), .CLK(clk_in), .RSTB(n7320), .Q(
        \FIFO[120][22] ) );
  DFFARX1 \FIFO_reg[120][21]  ( .D(n712), .CLK(clk_in), .RSTB(n7320), .Q(
        \FIFO[120][21] ) );
  DFFARX1 \FIFO_reg[120][20]  ( .D(n711), .CLK(clk_in), .RSTB(n7320), .Q(
        \FIFO[120][20] ) );
  DFFARX1 \FIFO_reg[120][19]  ( .D(n710), .CLK(clk_in), .RSTB(n7320), .Q(
        \FIFO[120][19] ) );
  DFFARX1 \FIFO_reg[120][18]  ( .D(n709), .CLK(clk_in), .RSTB(n7320), .Q(
        \FIFO[120][18] ) );
  DFFARX1 \FIFO_reg[120][17]  ( .D(n708), .CLK(clk_in), .RSTB(n7320), .Q(
        \FIFO[120][17] ) );
  DFFARX1 \FIFO_reg[120][16]  ( .D(n707), .CLK(clk_in), .RSTB(n7320), .Q(
        \FIFO[120][16] ) );
  DFFARX1 \FIFO_reg[120][15]  ( .D(n706), .CLK(clk_in), .RSTB(n7320), .Q(
        \FIFO[120][15] ) );
  DFFARX1 \FIFO_reg[120][14]  ( .D(n705), .CLK(clk_in), .RSTB(n7320), .Q(
        \FIFO[120][14] ) );
  DFFARX1 \FIFO_reg[120][13]  ( .D(n704), .CLK(clk_in), .RSTB(n7321), .Q(
        \FIFO[120][13] ) );
  DFFARX1 \FIFO_reg[120][12]  ( .D(n703), .CLK(clk_in), .RSTB(n7321), .Q(
        \FIFO[120][12] ) );
  DFFARX1 \FIFO_reg[120][11]  ( .D(n702), .CLK(clk_in), .RSTB(n7321), .Q(
        \FIFO[120][11] ) );
  DFFARX1 \FIFO_reg[120][10]  ( .D(n701), .CLK(clk_in), .RSTB(n7321), .Q(
        \FIFO[120][10] ) );
  DFFARX1 \FIFO_reg[120][9]  ( .D(n700), .CLK(clk_in), .RSTB(n7321), .Q(
        \FIFO[120][9] ) );
  DFFARX1 \FIFO_reg[120][8]  ( .D(n699), .CLK(clk_in), .RSTB(n7321), .Q(
        \FIFO[120][8] ) );
  DFFARX1 \FIFO_reg[120][7]  ( .D(n698), .CLK(clk_in), .RSTB(n7321), .Q(
        \FIFO[120][7] ) );
  DFFARX1 \FIFO_reg[120][6]  ( .D(n697), .CLK(clk_in), .RSTB(n7321), .Q(
        \FIFO[120][6] ) );
  DFFARX1 \FIFO_reg[120][5]  ( .D(n696), .CLK(clk_in), .RSTB(n7321), .Q(
        \FIFO[120][5] ) );
  DFFARX1 \FIFO_reg[120][4]  ( .D(n695), .CLK(clk_in), .RSTB(n7321), .Q(
        \FIFO[120][4] ) );
  DFFARX1 \FIFO_reg[120][3]  ( .D(n694), .CLK(clk_in), .RSTB(n7321), .Q(
        \FIFO[120][3] ) );
  DFFARX1 \FIFO_reg[120][2]  ( .D(n693), .CLK(clk_in), .RSTB(n7321), .Q(
        \FIFO[120][2] ) );
  DFFARX1 \FIFO_reg[120][1]  ( .D(n692), .CLK(clk_in), .RSTB(n7321), .Q(
        \FIFO[120][1] ) );
  DFFARX1 \FIFO_reg[120][0]  ( .D(n691), .CLK(clk_in), .RSTB(n7321), .Q(
        \FIFO[120][0] ) );
  DFFARX1 \FIFO_reg[121][31]  ( .D(n690), .CLK(clk_in), .RSTB(n7321), .Q(
        \FIFO[121][31] ) );
  DFFARX1 \FIFO_reg[121][30]  ( .D(n689), .CLK(clk_in), .RSTB(n7321), .Q(
        \FIFO[121][30] ) );
  DFFARX1 \FIFO_reg[121][29]  ( .D(n688), .CLK(clk_in), .RSTB(n7321), .Q(
        \FIFO[121][29] ) );
  DFFARX1 \FIFO_reg[121][28]  ( .D(n687), .CLK(clk_in), .RSTB(n7321), .Q(
        \FIFO[121][28] ) );
  DFFARX1 \FIFO_reg[121][27]  ( .D(n686), .CLK(clk_in), .RSTB(n7322), .Q(
        \FIFO[121][27] ) );
  DFFARX1 \FIFO_reg[121][26]  ( .D(n685), .CLK(clk_in), .RSTB(n7322), .Q(
        \FIFO[121][26] ) );
  DFFARX1 \FIFO_reg[121][25]  ( .D(n684), .CLK(clk_in), .RSTB(n7322), .Q(
        \FIFO[121][25] ) );
  DFFARX1 \FIFO_reg[121][24]  ( .D(n683), .CLK(clk_in), .RSTB(n7322), .Q(
        \FIFO[121][24] ) );
  DFFARX1 \FIFO_reg[121][23]  ( .D(n682), .CLK(clk_in), .RSTB(n7322), .Q(
        \FIFO[121][23] ) );
  DFFARX1 \FIFO_reg[121][22]  ( .D(n681), .CLK(clk_in), .RSTB(n7322), .Q(
        \FIFO[121][22] ) );
  DFFARX1 \FIFO_reg[121][21]  ( .D(n680), .CLK(clk_in), .RSTB(n7322), .Q(
        \FIFO[121][21] ) );
  DFFARX1 \FIFO_reg[121][20]  ( .D(n679), .CLK(clk_in), .RSTB(n7322), .Q(
        \FIFO[121][20] ) );
  DFFARX1 \FIFO_reg[121][19]  ( .D(n678), .CLK(clk_in), .RSTB(n7322), .Q(
        \FIFO[121][19] ) );
  DFFARX1 \FIFO_reg[121][18]  ( .D(n677), .CLK(clk_in), .RSTB(n7322), .Q(
        \FIFO[121][18] ) );
  DFFARX1 \FIFO_reg[121][17]  ( .D(n676), .CLK(clk_in), .RSTB(n7322), .Q(
        \FIFO[121][17] ) );
  DFFARX1 \FIFO_reg[121][16]  ( .D(n675), .CLK(clk_in), .RSTB(n7322), .Q(
        \FIFO[121][16] ) );
  DFFARX1 \FIFO_reg[121][15]  ( .D(n674), .CLK(clk_in), .RSTB(n7322), .Q(
        \FIFO[121][15] ) );
  DFFARX1 \FIFO_reg[121][14]  ( .D(n673), .CLK(clk_in), .RSTB(n7322), .Q(
        \FIFO[121][14] ) );
  DFFARX1 \FIFO_reg[121][13]  ( .D(n672), .CLK(clk_in), .RSTB(n7322), .Q(
        \FIFO[121][13] ) );
  DFFARX1 \FIFO_reg[121][12]  ( .D(n671), .CLK(clk_in), .RSTB(n7322), .Q(
        \FIFO[121][12] ) );
  DFFARX1 \FIFO_reg[121][11]  ( .D(n670), .CLK(clk_in), .RSTB(n7322), .Q(
        \FIFO[121][11] ) );
  DFFARX1 \FIFO_reg[121][10]  ( .D(n669), .CLK(clk_in), .RSTB(n7322), .Q(
        \FIFO[121][10] ) );
  DFFARX1 \FIFO_reg[121][9]  ( .D(n668), .CLK(clk_in), .RSTB(n7323), .Q(
        \FIFO[121][9] ) );
  DFFARX1 \FIFO_reg[121][8]  ( .D(n667), .CLK(clk_in), .RSTB(n7323), .Q(
        \FIFO[121][8] ) );
  DFFARX1 \FIFO_reg[121][7]  ( .D(n666), .CLK(clk_in), .RSTB(n7323), .Q(
        \FIFO[121][7] ) );
  DFFARX1 \FIFO_reg[121][6]  ( .D(n665), .CLK(clk_in), .RSTB(n7323), .Q(
        \FIFO[121][6] ) );
  DFFARX1 \FIFO_reg[121][5]  ( .D(n664), .CLK(clk_in), .RSTB(n7323), .Q(
        \FIFO[121][5] ) );
  DFFARX1 \FIFO_reg[121][4]  ( .D(n663), .CLK(clk_in), .RSTB(n7323), .Q(
        \FIFO[121][4] ) );
  DFFARX1 \FIFO_reg[121][3]  ( .D(n662), .CLK(clk_in), .RSTB(n7323), .Q(
        \FIFO[121][3] ) );
  DFFARX1 \FIFO_reg[121][2]  ( .D(n661), .CLK(clk_in), .RSTB(n7323), .Q(
        \FIFO[121][2] ) );
  DFFARX1 \FIFO_reg[121][1]  ( .D(n660), .CLK(clk_in), .RSTB(n7323), .Q(
        \FIFO[121][1] ) );
  DFFARX1 \FIFO_reg[121][0]  ( .D(n659), .CLK(clk_in), .RSTB(n7323), .Q(
        \FIFO[121][0] ) );
  DFFARX1 \FIFO_reg[122][31]  ( .D(n658), .CLK(clk_in), .RSTB(n7323), .Q(
        \FIFO[122][31] ) );
  DFFARX1 \FIFO_reg[122][30]  ( .D(n657), .CLK(clk_in), .RSTB(n7323), .Q(
        \FIFO[122][30] ) );
  DFFARX1 \FIFO_reg[122][29]  ( .D(n656), .CLK(clk_in), .RSTB(n7323), .Q(
        \FIFO[122][29] ) );
  DFFARX1 \FIFO_reg[122][28]  ( .D(n655), .CLK(clk_in), .RSTB(n7323), .Q(
        \FIFO[122][28] ) );
  DFFARX1 \FIFO_reg[122][27]  ( .D(n654), .CLK(clk_in), .RSTB(n7323), .Q(
        \FIFO[122][27] ) );
  DFFARX1 \FIFO_reg[122][26]  ( .D(n653), .CLK(clk_in), .RSTB(n7323), .Q(
        \FIFO[122][26] ) );
  DFFARX1 \FIFO_reg[122][25]  ( .D(n652), .CLK(clk_in), .RSTB(n7323), .Q(
        \FIFO[122][25] ) );
  DFFARX1 \FIFO_reg[122][24]  ( .D(n651), .CLK(clk_in), .RSTB(n7323), .Q(
        \FIFO[122][24] ) );
  DFFARX1 \FIFO_reg[122][23]  ( .D(n650), .CLK(clk_in), .RSTB(n7324), .Q(
        \FIFO[122][23] ) );
  DFFARX1 \FIFO_reg[122][22]  ( .D(n649), .CLK(clk_in), .RSTB(n7324), .Q(
        \FIFO[122][22] ) );
  DFFARX1 \FIFO_reg[122][21]  ( .D(n648), .CLK(clk_in), .RSTB(n7324), .Q(
        \FIFO[122][21] ) );
  DFFARX1 \FIFO_reg[122][20]  ( .D(n647), .CLK(clk_in), .RSTB(n7324), .Q(
        \FIFO[122][20] ) );
  DFFARX1 \FIFO_reg[122][19]  ( .D(n646), .CLK(clk_in), .RSTB(n7324), .Q(
        \FIFO[122][19] ) );
  DFFARX1 \FIFO_reg[122][18]  ( .D(n645), .CLK(clk_in), .RSTB(n7324), .Q(
        \FIFO[122][18] ) );
  DFFARX1 \FIFO_reg[122][17]  ( .D(n644), .CLK(clk_in), .RSTB(n7324), .Q(
        \FIFO[122][17] ) );
  DFFARX1 \FIFO_reg[122][16]  ( .D(n643), .CLK(clk_in), .RSTB(n7324), .Q(
        \FIFO[122][16] ) );
  DFFARX1 \FIFO_reg[122][15]  ( .D(n642), .CLK(clk_in), .RSTB(n7324), .Q(
        \FIFO[122][15] ) );
  DFFARX1 \FIFO_reg[122][14]  ( .D(n641), .CLK(clk_in), .RSTB(n7324), .Q(
        \FIFO[122][14] ) );
  DFFARX1 \FIFO_reg[122][13]  ( .D(n640), .CLK(clk_in), .RSTB(n7324), .Q(
        \FIFO[122][13] ) );
  DFFARX1 \FIFO_reg[122][12]  ( .D(n639), .CLK(clk_in), .RSTB(n7324), .Q(
        \FIFO[122][12] ) );
  DFFARX1 \FIFO_reg[122][11]  ( .D(n638), .CLK(clk_in), .RSTB(n7324), .Q(
        \FIFO[122][11] ) );
  DFFARX1 \FIFO_reg[122][10]  ( .D(n637), .CLK(clk_in), .RSTB(n7324), .Q(
        \FIFO[122][10] ) );
  DFFARX1 \FIFO_reg[122][9]  ( .D(n636), .CLK(clk_in), .RSTB(n7324), .Q(
        \FIFO[122][9] ) );
  DFFARX1 \FIFO_reg[122][8]  ( .D(n635), .CLK(clk_in), .RSTB(n7324), .Q(
        \FIFO[122][8] ) );
  DFFARX1 \FIFO_reg[122][7]  ( .D(n634), .CLK(clk_in), .RSTB(n7324), .Q(
        \FIFO[122][7] ) );
  DFFARX1 \FIFO_reg[122][6]  ( .D(n633), .CLK(clk_in), .RSTB(n7324), .Q(
        \FIFO[122][6] ) );
  DFFARX1 \FIFO_reg[122][5]  ( .D(n632), .CLK(clk_in), .RSTB(n7325), .Q(
        \FIFO[122][5] ) );
  DFFARX1 \FIFO_reg[122][4]  ( .D(n631), .CLK(clk_in), .RSTB(n7325), .Q(
        \FIFO[122][4] ) );
  DFFARX1 \FIFO_reg[122][3]  ( .D(n630), .CLK(clk_in), .RSTB(n7325), .Q(
        \FIFO[122][3] ) );
  DFFARX1 \FIFO_reg[122][2]  ( .D(n629), .CLK(clk_in), .RSTB(n7325), .Q(
        \FIFO[122][2] ) );
  DFFARX1 \FIFO_reg[122][1]  ( .D(n628), .CLK(clk_in), .RSTB(n7325), .Q(
        \FIFO[122][1] ) );
  DFFARX1 \FIFO_reg[122][0]  ( .D(n627), .CLK(clk_in), .RSTB(n7325), .Q(
        \FIFO[122][0] ) );
  DFFARX1 \FIFO_reg[123][31]  ( .D(n626), .CLK(clk_in), .RSTB(n7325), .Q(
        \FIFO[123][31] ) );
  DFFARX1 \FIFO_reg[123][30]  ( .D(n625), .CLK(clk_in), .RSTB(n7325), .Q(
        \FIFO[123][30] ) );
  DFFARX1 \FIFO_reg[123][29]  ( .D(n624), .CLK(clk_in), .RSTB(n7325), .Q(
        \FIFO[123][29] ) );
  DFFARX1 \FIFO_reg[123][28]  ( .D(n623), .CLK(clk_in), .RSTB(n7325), .Q(
        \FIFO[123][28] ) );
  DFFARX1 \FIFO_reg[123][27]  ( .D(n622), .CLK(clk_in), .RSTB(n7325), .Q(
        \FIFO[123][27] ) );
  DFFARX1 \FIFO_reg[123][26]  ( .D(n621), .CLK(clk_in), .RSTB(n7325), .Q(
        \FIFO[123][26] ) );
  DFFARX1 \FIFO_reg[123][25]  ( .D(n620), .CLK(clk_in), .RSTB(n7325), .Q(
        \FIFO[123][25] ) );
  DFFARX1 \FIFO_reg[123][24]  ( .D(n619), .CLK(clk_in), .RSTB(n7325), .Q(
        \FIFO[123][24] ) );
  DFFARX1 \FIFO_reg[123][23]  ( .D(n618), .CLK(clk_in), .RSTB(n7325), .Q(
        \FIFO[123][23] ) );
  DFFARX1 \FIFO_reg[123][22]  ( .D(n617), .CLK(clk_in), .RSTB(n7325), .Q(
        \FIFO[123][22] ) );
  DFFARX1 \FIFO_reg[123][21]  ( .D(n616), .CLK(clk_in), .RSTB(n7325), .Q(
        \FIFO[123][21] ) );
  DFFARX1 \FIFO_reg[123][20]  ( .D(n615), .CLK(clk_in), .RSTB(n7325), .Q(
        \FIFO[123][20] ) );
  DFFARX1 \FIFO_reg[123][19]  ( .D(n614), .CLK(clk_in), .RSTB(n7326), .Q(
        \FIFO[123][19] ) );
  DFFARX1 \FIFO_reg[123][18]  ( .D(n613), .CLK(clk_in), .RSTB(n7326), .Q(
        \FIFO[123][18] ) );
  DFFARX1 \FIFO_reg[123][17]  ( .D(n612), .CLK(clk_in), .RSTB(n7326), .Q(
        \FIFO[123][17] ) );
  DFFARX1 \FIFO_reg[123][16]  ( .D(n611), .CLK(clk_in), .RSTB(n7326), .Q(
        \FIFO[123][16] ) );
  DFFARX1 \FIFO_reg[123][15]  ( .D(n610), .CLK(clk_in), .RSTB(n7326), .Q(
        \FIFO[123][15] ) );
  DFFARX1 \FIFO_reg[123][14]  ( .D(n609), .CLK(clk_in), .RSTB(n7326), .Q(
        \FIFO[123][14] ) );
  DFFARX1 \FIFO_reg[123][13]  ( .D(n608), .CLK(clk_in), .RSTB(n7326), .Q(
        \FIFO[123][13] ) );
  DFFARX1 \FIFO_reg[123][12]  ( .D(n607), .CLK(clk_in), .RSTB(n7326), .Q(
        \FIFO[123][12] ) );
  DFFARX1 \FIFO_reg[123][11]  ( .D(n606), .CLK(clk_in), .RSTB(n7326), .Q(
        \FIFO[123][11] ) );
  DFFARX1 \FIFO_reg[123][10]  ( .D(n605), .CLK(clk_in), .RSTB(n7326), .Q(
        \FIFO[123][10] ) );
  DFFARX1 \FIFO_reg[123][9]  ( .D(n604), .CLK(clk_in), .RSTB(n7326), .Q(
        \FIFO[123][9] ) );
  DFFARX1 \FIFO_reg[123][8]  ( .D(n603), .CLK(clk_in), .RSTB(n7326), .Q(
        \FIFO[123][8] ) );
  DFFARX1 \FIFO_reg[123][7]  ( .D(n602), .CLK(clk_in), .RSTB(n7326), .Q(
        \FIFO[123][7] ) );
  DFFARX1 \FIFO_reg[123][6]  ( .D(n601), .CLK(clk_in), .RSTB(n7326), .Q(
        \FIFO[123][6] ) );
  DFFARX1 \FIFO_reg[123][5]  ( .D(n600), .CLK(clk_in), .RSTB(n7326), .Q(
        \FIFO[123][5] ) );
  DFFARX1 \FIFO_reg[123][4]  ( .D(n599), .CLK(clk_in), .RSTB(n7326), .Q(
        \FIFO[123][4] ) );
  DFFARX1 \FIFO_reg[123][3]  ( .D(n598), .CLK(clk_in), .RSTB(n7326), .Q(
        \FIFO[123][3] ) );
  DFFARX1 \FIFO_reg[123][2]  ( .D(n597), .CLK(clk_in), .RSTB(n7326), .Q(
        \FIFO[123][2] ) );
  DFFARX1 \FIFO_reg[123][1]  ( .D(n596), .CLK(clk_in), .RSTB(n7327), .Q(
        \FIFO[123][1] ) );
  DFFARX1 \FIFO_reg[123][0]  ( .D(n595), .CLK(clk_in), .RSTB(n7327), .Q(
        \FIFO[123][0] ) );
  DFFARX1 \FIFO_reg[124][31]  ( .D(n594), .CLK(clk_in), .RSTB(n7327), .Q(
        \FIFO[124][31] ) );
  DFFARX1 \FIFO_reg[124][30]  ( .D(n593), .CLK(clk_in), .RSTB(n7327), .Q(
        \FIFO[124][30] ) );
  DFFARX1 \FIFO_reg[124][29]  ( .D(n592), .CLK(clk_in), .RSTB(n7327), .Q(
        \FIFO[124][29] ) );
  DFFARX1 \FIFO_reg[124][28]  ( .D(n591), .CLK(clk_in), .RSTB(n7327), .Q(
        \FIFO[124][28] ) );
  DFFARX1 \FIFO_reg[124][27]  ( .D(n590), .CLK(clk_in), .RSTB(n7327), .Q(
        \FIFO[124][27] ) );
  DFFARX1 \FIFO_reg[124][26]  ( .D(n589), .CLK(clk_in), .RSTB(n7327), .Q(
        \FIFO[124][26] ) );
  DFFARX1 \FIFO_reg[124][25]  ( .D(n588), .CLK(clk_in), .RSTB(n7327), .Q(
        \FIFO[124][25] ) );
  DFFARX1 \FIFO_reg[124][24]  ( .D(n587), .CLK(clk_in), .RSTB(n7327), .Q(
        \FIFO[124][24] ) );
  DFFARX1 \FIFO_reg[124][23]  ( .D(n586), .CLK(clk_in), .RSTB(n7327), .Q(
        \FIFO[124][23] ) );
  DFFARX1 \FIFO_reg[124][22]  ( .D(n585), .CLK(clk_in), .RSTB(n7327), .Q(
        \FIFO[124][22] ) );
  DFFARX1 \FIFO_reg[124][21]  ( .D(n584), .CLK(clk_in), .RSTB(n7327), .Q(
        \FIFO[124][21] ) );
  DFFARX1 \FIFO_reg[124][20]  ( .D(n583), .CLK(clk_in), .RSTB(n7327), .Q(
        \FIFO[124][20] ) );
  DFFARX1 \FIFO_reg[124][19]  ( .D(n582), .CLK(clk_in), .RSTB(n7327), .Q(
        \FIFO[124][19] ) );
  DFFARX1 \FIFO_reg[124][18]  ( .D(n581), .CLK(clk_in), .RSTB(n7327), .Q(
        \FIFO[124][18] ) );
  DFFARX1 \FIFO_reg[124][17]  ( .D(n580), .CLK(clk_in), .RSTB(n7327), .Q(
        \FIFO[124][17] ) );
  DFFARX1 \FIFO_reg[124][16]  ( .D(n579), .CLK(clk_in), .RSTB(n7327), .Q(
        \FIFO[124][16] ) );
  DFFARX1 \FIFO_reg[124][15]  ( .D(n578), .CLK(clk_in), .RSTB(n7328), .Q(
        \FIFO[124][15] ) );
  DFFARX1 \FIFO_reg[124][14]  ( .D(n577), .CLK(clk_in), .RSTB(n7328), .Q(
        \FIFO[124][14] ) );
  DFFARX1 \FIFO_reg[124][13]  ( .D(n576), .CLK(clk_in), .RSTB(n7328), .Q(
        \FIFO[124][13] ) );
  DFFARX1 \FIFO_reg[124][12]  ( .D(n575), .CLK(clk_in), .RSTB(n7328), .Q(
        \FIFO[124][12] ) );
  DFFARX1 \FIFO_reg[124][11]  ( .D(n574), .CLK(clk_in), .RSTB(n7328), .Q(
        \FIFO[124][11] ) );
  DFFARX1 \FIFO_reg[124][10]  ( .D(n573), .CLK(clk_in), .RSTB(n7328), .Q(
        \FIFO[124][10] ) );
  DFFARX1 \FIFO_reg[124][9]  ( .D(n572), .CLK(clk_in), .RSTB(n7328), .Q(
        \FIFO[124][9] ) );
  DFFARX1 \FIFO_reg[124][8]  ( .D(n571), .CLK(clk_in), .RSTB(n7328), .Q(
        \FIFO[124][8] ) );
  DFFARX1 \FIFO_reg[124][7]  ( .D(n570), .CLK(clk_in), .RSTB(n7328), .Q(
        \FIFO[124][7] ) );
  DFFARX1 \FIFO_reg[124][6]  ( .D(n569), .CLK(clk_in), .RSTB(n7328), .Q(
        \FIFO[124][6] ) );
  DFFARX1 \FIFO_reg[124][5]  ( .D(n568), .CLK(clk_in), .RSTB(n7328), .Q(
        \FIFO[124][5] ) );
  DFFARX1 \FIFO_reg[124][4]  ( .D(n567), .CLK(clk_in), .RSTB(n7328), .Q(
        \FIFO[124][4] ) );
  DFFARX1 \FIFO_reg[124][3]  ( .D(n566), .CLK(clk_in), .RSTB(n7328), .Q(
        \FIFO[124][3] ) );
  DFFARX1 \FIFO_reg[124][2]  ( .D(n565), .CLK(clk_in), .RSTB(n7328), .Q(
        \FIFO[124][2] ) );
  DFFARX1 \FIFO_reg[124][1]  ( .D(n564), .CLK(clk_in), .RSTB(n7328), .Q(
        \FIFO[124][1] ) );
  DFFARX1 \FIFO_reg[124][0]  ( .D(n563), .CLK(clk_in), .RSTB(n7328), .Q(
        \FIFO[124][0] ) );
  DFFARX1 \FIFO_reg[125][31]  ( .D(n562), .CLK(clk_in), .RSTB(n7328), .Q(
        \FIFO[125][31] ) );
  DFFARX1 \FIFO_reg[125][30]  ( .D(n561), .CLK(clk_in), .RSTB(n7328), .Q(
        \FIFO[125][30] ) );
  DFFARX1 \FIFO_reg[125][29]  ( .D(n560), .CLK(clk_in), .RSTB(n7329), .Q(
        \FIFO[125][29] ) );
  DFFARX1 \FIFO_reg[125][28]  ( .D(n559), .CLK(clk_in), .RSTB(n7329), .Q(
        \FIFO[125][28] ) );
  DFFARX1 \FIFO_reg[125][27]  ( .D(n558), .CLK(clk_in), .RSTB(n7329), .Q(
        \FIFO[125][27] ) );
  DFFARX1 \FIFO_reg[125][26]  ( .D(n557), .CLK(clk_in), .RSTB(n7329), .Q(
        \FIFO[125][26] ) );
  DFFARX1 \FIFO_reg[125][25]  ( .D(n556), .CLK(clk_in), .RSTB(n7329), .Q(
        \FIFO[125][25] ) );
  DFFARX1 \FIFO_reg[125][24]  ( .D(n555), .CLK(clk_in), .RSTB(n7329), .Q(
        \FIFO[125][24] ) );
  DFFARX1 \FIFO_reg[125][23]  ( .D(n554), .CLK(clk_in), .RSTB(n7329), .Q(
        \FIFO[125][23] ) );
  DFFARX1 \FIFO_reg[125][22]  ( .D(n553), .CLK(clk_in), .RSTB(n7329), .Q(
        \FIFO[125][22] ) );
  DFFARX1 \FIFO_reg[125][21]  ( .D(n552), .CLK(clk_in), .RSTB(n7329), .Q(
        \FIFO[125][21] ) );
  DFFARX1 \FIFO_reg[125][20]  ( .D(n551), .CLK(clk_in), .RSTB(n7329), .Q(
        \FIFO[125][20] ) );
  DFFARX1 \FIFO_reg[125][19]  ( .D(n550), .CLK(clk_in), .RSTB(n7329), .Q(
        \FIFO[125][19] ) );
  DFFARX1 \FIFO_reg[125][18]  ( .D(n549), .CLK(clk_in), .RSTB(n7329), .Q(
        \FIFO[125][18] ) );
  DFFARX1 \FIFO_reg[125][17]  ( .D(n548), .CLK(clk_in), .RSTB(n7329), .Q(
        \FIFO[125][17] ) );
  DFFARX1 \FIFO_reg[125][16]  ( .D(n547), .CLK(clk_in), .RSTB(n7329), .Q(
        \FIFO[125][16] ) );
  DFFARX1 \FIFO_reg[125][15]  ( .D(n546), .CLK(clk_in), .RSTB(n7329), .Q(
        \FIFO[125][15] ) );
  DFFARX1 \FIFO_reg[125][14]  ( .D(n545), .CLK(clk_in), .RSTB(n7329), .Q(
        \FIFO[125][14] ) );
  DFFARX1 \FIFO_reg[125][13]  ( .D(n544), .CLK(clk_in), .RSTB(n7329), .Q(
        \FIFO[125][13] ) );
  DFFARX1 \FIFO_reg[125][12]  ( .D(n543), .CLK(clk_in), .RSTB(n7329), .Q(
        \FIFO[125][12] ) );
  DFFARX1 \FIFO_reg[125][11]  ( .D(n542), .CLK(clk_in), .RSTB(n7330), .Q(
        \FIFO[125][11] ) );
  DFFARX1 \FIFO_reg[125][10]  ( .D(n541), .CLK(clk_in), .RSTB(n7330), .Q(
        \FIFO[125][10] ) );
  DFFARX1 \FIFO_reg[125][9]  ( .D(n540), .CLK(clk_in), .RSTB(n7330), .Q(
        \FIFO[125][9] ) );
  DFFARX1 \FIFO_reg[125][8]  ( .D(n539), .CLK(clk_in), .RSTB(n7330), .Q(
        \FIFO[125][8] ) );
  DFFARX1 \FIFO_reg[125][7]  ( .D(n538), .CLK(clk_in), .RSTB(n7330), .Q(
        \FIFO[125][7] ) );
  DFFARX1 \FIFO_reg[125][6]  ( .D(n537), .CLK(clk_in), .RSTB(n7330), .Q(
        \FIFO[125][6] ) );
  DFFARX1 \FIFO_reg[125][5]  ( .D(n536), .CLK(clk_in), .RSTB(n7330), .Q(
        \FIFO[125][5] ) );
  DFFARX1 \FIFO_reg[125][4]  ( .D(n535), .CLK(clk_in), .RSTB(n7330), .Q(
        \FIFO[125][4] ) );
  DFFARX1 \FIFO_reg[125][3]  ( .D(n534), .CLK(clk_in), .RSTB(n7330), .Q(
        \FIFO[125][3] ) );
  DFFARX1 \FIFO_reg[125][2]  ( .D(n533), .CLK(clk_in), .RSTB(n7330), .Q(
        \FIFO[125][2] ) );
  DFFARX1 \FIFO_reg[125][1]  ( .D(n532), .CLK(clk_in), .RSTB(n7330), .Q(
        \FIFO[125][1] ) );
  DFFARX1 \FIFO_reg[125][0]  ( .D(n531), .CLK(clk_in), .RSTB(n7330), .Q(
        \FIFO[125][0] ) );
  DFFARX1 \FIFO_reg[126][31]  ( .D(n530), .CLK(clk_in), .RSTB(n7330), .Q(
        \FIFO[126][31] ) );
  DFFARX1 \FIFO_reg[126][30]  ( .D(n529), .CLK(clk_in), .RSTB(n7330), .Q(
        \FIFO[126][30] ) );
  DFFARX1 \FIFO_reg[126][29]  ( .D(n528), .CLK(clk_in), .RSTB(n7330), .Q(
        \FIFO[126][29] ) );
  DFFARX1 \FIFO_reg[126][28]  ( .D(n527), .CLK(clk_in), .RSTB(n7330), .Q(
        \FIFO[126][28] ) );
  DFFARX1 \FIFO_reg[126][27]  ( .D(n526), .CLK(clk_in), .RSTB(n7330), .Q(
        \FIFO[126][27] ) );
  DFFARX1 \FIFO_reg[126][26]  ( .D(n525), .CLK(clk_in), .RSTB(n7330), .Q(
        \FIFO[126][26] ) );
  DFFARX1 \FIFO_reg[126][25]  ( .D(n524), .CLK(clk_in), .RSTB(n7331), .Q(
        \FIFO[126][25] ) );
  DFFARX1 \FIFO_reg[126][24]  ( .D(n523), .CLK(clk_in), .RSTB(n7331), .Q(
        \FIFO[126][24] ) );
  DFFARX1 \FIFO_reg[126][23]  ( .D(n522), .CLK(clk_in), .RSTB(n7331), .Q(
        \FIFO[126][23] ) );
  DFFARX1 \FIFO_reg[126][22]  ( .D(n521), .CLK(clk_in), .RSTB(n7331), .Q(
        \FIFO[126][22] ) );
  DFFARX1 \FIFO_reg[126][21]  ( .D(n520), .CLK(clk_in), .RSTB(n7331), .Q(
        \FIFO[126][21] ) );
  DFFARX1 \FIFO_reg[126][20]  ( .D(n519), .CLK(clk_in), .RSTB(n7331), .Q(
        \FIFO[126][20] ) );
  DFFARX1 \FIFO_reg[126][19]  ( .D(n518), .CLK(clk_in), .RSTB(n7331), .Q(
        \FIFO[126][19] ) );
  DFFARX1 \FIFO_reg[126][18]  ( .D(n517), .CLK(clk_in), .RSTB(n7331), .Q(
        \FIFO[126][18] ) );
  DFFARX1 \FIFO_reg[126][17]  ( .D(n516), .CLK(clk_in), .RSTB(n7331), .Q(
        \FIFO[126][17] ) );
  DFFARX1 \FIFO_reg[126][16]  ( .D(n515), .CLK(clk_in), .RSTB(n7331), .Q(
        \FIFO[126][16] ) );
  DFFARX1 \FIFO_reg[126][15]  ( .D(n514), .CLK(clk_in), .RSTB(n7331), .Q(
        \FIFO[126][15] ) );
  DFFARX1 \FIFO_reg[126][14]  ( .D(n513), .CLK(clk_in), .RSTB(n7331), .Q(
        \FIFO[126][14] ) );
  DFFARX1 \FIFO_reg[126][13]  ( .D(n512), .CLK(clk_in), .RSTB(n7331), .Q(
        \FIFO[126][13] ) );
  DFFARX1 \FIFO_reg[126][12]  ( .D(n511), .CLK(clk_in), .RSTB(n7331), .Q(
        \FIFO[126][12] ) );
  DFFARX1 \FIFO_reg[126][11]  ( .D(n510), .CLK(clk_in), .RSTB(n7331), .Q(
        \FIFO[126][11] ) );
  DFFARX1 \FIFO_reg[126][10]  ( .D(n509), .CLK(clk_in), .RSTB(n7331), .Q(
        \FIFO[126][10] ) );
  DFFARX1 \FIFO_reg[126][9]  ( .D(n508), .CLK(clk_in), .RSTB(n7331), .Q(
        \FIFO[126][9] ) );
  DFFARX1 \FIFO_reg[126][8]  ( .D(n507), .CLK(clk_in), .RSTB(n7331), .Q(
        \FIFO[126][8] ) );
  DFFARX1 \FIFO_reg[126][7]  ( .D(n506), .CLK(clk_in), .RSTB(n7332), .Q(
        \FIFO[126][7] ) );
  DFFARX1 \FIFO_reg[126][6]  ( .D(n505), .CLK(clk_in), .RSTB(n7332), .Q(
        \FIFO[126][6] ) );
  DFFARX1 \FIFO_reg[126][5]  ( .D(n504), .CLK(clk_in), .RSTB(n7332), .Q(
        \FIFO[126][5] ) );
  DFFARX1 \FIFO_reg[126][4]  ( .D(n503), .CLK(clk_in), .RSTB(n7332), .Q(
        \FIFO[126][4] ) );
  DFFARX1 \FIFO_reg[126][3]  ( .D(n502), .CLK(clk_in), .RSTB(n7332), .Q(
        \FIFO[126][3] ) );
  DFFARX1 \FIFO_reg[126][2]  ( .D(n501), .CLK(clk_in), .RSTB(n7332), .Q(
        \FIFO[126][2] ) );
  DFFARX1 \FIFO_reg[126][1]  ( .D(n500), .CLK(clk_in), .RSTB(n7332), .Q(
        \FIFO[126][1] ) );
  DFFARX1 \FIFO_reg[126][0]  ( .D(n499), .CLK(clk_in), .RSTB(n7332), .Q(
        \FIFO[126][0] ) );
  DFFARX1 \FIFO_reg[127][31]  ( .D(n498), .CLK(clk_in), .RSTB(n7332), .Q(
        \FIFO[127][31] ) );
  DFFARX1 \FIFO_reg[127][30]  ( .D(n497), .CLK(clk_in), .RSTB(n7332), .Q(
        \FIFO[127][30] ) );
  DFFARX1 \FIFO_reg[127][29]  ( .D(n496), .CLK(clk_in), .RSTB(n7332), .Q(
        \FIFO[127][29] ) );
  DFFARX1 \FIFO_reg[127][28]  ( .D(n495), .CLK(clk_in), .RSTB(n7332), .Q(
        \FIFO[127][28] ) );
  DFFARX1 \FIFO_reg[127][27]  ( .D(n494), .CLK(clk_in), .RSTB(n7332), .Q(
        \FIFO[127][27] ) );
  DFFARX1 \FIFO_reg[127][26]  ( .D(n493), .CLK(clk_in), .RSTB(n7332), .Q(
        \FIFO[127][26] ) );
  DFFARX1 \FIFO_reg[127][25]  ( .D(n492), .CLK(clk_in), .RSTB(n7332), .Q(
        \FIFO[127][25] ) );
  DFFARX1 \FIFO_reg[127][24]  ( .D(n491), .CLK(clk_in), .RSTB(n7332), .Q(
        \FIFO[127][24] ) );
  DFFARX1 \FIFO_reg[127][23]  ( .D(n490), .CLK(clk_in), .RSTB(n7332), .Q(
        \FIFO[127][23] ) );
  DFFARX1 \FIFO_reg[127][22]  ( .D(n489), .CLK(clk_in), .RSTB(n7332), .Q(
        \FIFO[127][22] ) );
  DFFARX1 \FIFO_reg[127][21]  ( .D(n488), .CLK(clk_in), .RSTB(n7333), .Q(
        \FIFO[127][21] ) );
  DFFARX1 \FIFO_reg[127][20]  ( .D(n487), .CLK(clk_in), .RSTB(n7333), .Q(
        \FIFO[127][20] ) );
  DFFARX1 \FIFO_reg[127][19]  ( .D(n486), .CLK(clk_in), .RSTB(n7333), .Q(
        \FIFO[127][19] ) );
  DFFARX1 \FIFO_reg[127][18]  ( .D(n485), .CLK(clk_in), .RSTB(n7333), .Q(
        \FIFO[127][18] ) );
  DFFARX1 \FIFO_reg[127][17]  ( .D(n484), .CLK(clk_in), .RSTB(n7333), .Q(
        \FIFO[127][17] ) );
  DFFARX1 \FIFO_reg[127][16]  ( .D(n483), .CLK(clk_in), .RSTB(n7333), .Q(
        \FIFO[127][16] ) );
  DFFARX1 \FIFO_reg[127][15]  ( .D(n482), .CLK(clk_in), .RSTB(n7333), .Q(
        \FIFO[127][15] ) );
  DFFARX1 \FIFO_reg[127][14]  ( .D(n481), .CLK(clk_in), .RSTB(n7333), .Q(
        \FIFO[127][14] ) );
  DFFARX1 \FIFO_reg[127][13]  ( .D(n480), .CLK(clk_in), .RSTB(n7333), .Q(
        \FIFO[127][13] ) );
  DFFARX1 \FIFO_reg[127][12]  ( .D(n479), .CLK(clk_in), .RSTB(n7333), .Q(
        \FIFO[127][12] ) );
  DFFARX1 \FIFO_reg[127][11]  ( .D(n478), .CLK(clk_in), .RSTB(n7333), .Q(
        \FIFO[127][11] ) );
  DFFARX1 \FIFO_reg[127][10]  ( .D(n477), .CLK(clk_in), .RSTB(n7333), .Q(
        \FIFO[127][10] ) );
  DFFARX1 \FIFO_reg[127][9]  ( .D(n476), .CLK(clk_in), .RSTB(n7333), .Q(
        \FIFO[127][9] ) );
  DFFARX1 \FIFO_reg[127][8]  ( .D(n475), .CLK(clk_in), .RSTB(n7333), .Q(
        \FIFO[127][8] ) );
  DFFARX1 \FIFO_reg[127][7]  ( .D(n474), .CLK(clk_in), .RSTB(n7333), .Q(
        \FIFO[127][7] ) );
  DFFARX1 \FIFO_reg[127][6]  ( .D(n473), .CLK(clk_in), .RSTB(n7333), .Q(
        \FIFO[127][6] ) );
  DFFARX1 \FIFO_reg[127][5]  ( .D(n472), .CLK(clk_in), .RSTB(n7333), .Q(
        \FIFO[127][5] ) );
  DFFARX1 \FIFO_reg[127][4]  ( .D(n471), .CLK(clk_in), .RSTB(n7333), .Q(
        \FIFO[127][4] ) );
  DFFARX1 \FIFO_reg[127][3]  ( .D(n470), .CLK(clk_in), .RSTB(rst), .Q(
        \FIFO[127][3] ) );
  DFFARX1 \FIFO_reg[127][2]  ( .D(n469), .CLK(clk_in), .RSTB(rst), .Q(
        \FIFO[127][2] ) );
  DFFARX1 \FIFO_reg[127][1]  ( .D(n468), .CLK(clk_in), .RSTB(rst), .Q(
        \FIFO[127][1] ) );
  DFFARX1 \FIFO_reg[127][0]  ( .D(n467), .CLK(clk_in), .RSTB(rst), .Q(
        \FIFO[127][0] ) );
  DFFASRX1 \dataOut_reg[31]  ( .D(n464), .CLK(clk_out), .RSTB(n85), .SETB(n117), .Q(dataOut[31]) );
  DFFASRX1 \dataOut_reg[30]  ( .D(N283), .CLK(clk_out), .RSTB(n84), .SETB(n116), .Q(dataOut[30]) );
  DFFASRX1 \dataOut_reg[29]  ( .D(N282), .CLK(clk_out), .RSTB(n83), .SETB(n115), .Q(dataOut[29]) );
  DFFASRX1 \dataOut_reg[28]  ( .D(N281), .CLK(clk_out), .RSTB(n82), .SETB(n114), .Q(dataOut[28]) );
  DFFASRX1 \dataOut_reg[27]  ( .D(N280), .CLK(clk_out), .RSTB(n81), .SETB(n113), .Q(dataOut[27]) );
  DFFASRX1 \dataOut_reg[26]  ( .D(N279), .CLK(clk_out), .RSTB(n80), .SETB(n112), .Q(dataOut[26]) );
  DFFASRX1 \dataOut_reg[25]  ( .D(N278), .CLK(clk_out), .RSTB(n79), .SETB(n111), .Q(dataOut[25]) );
  DFFASRX1 \dataOut_reg[24]  ( .D(N277), .CLK(clk_out), .RSTB(n78), .SETB(n110), .Q(dataOut[24]) );
  DFFASRX1 \dataOut_reg[23]  ( .D(N276), .CLK(clk_out), .RSTB(n77), .SETB(n109), .Q(dataOut[23]) );
  DFFASRX1 \dataOut_reg[22]  ( .D(N275), .CLK(clk_out), .RSTB(n76), .SETB(n108), .Q(dataOut[22]) );
  DFFASRX1 \dataOut_reg[21]  ( .D(N274), .CLK(clk_out), .RSTB(n75), .SETB(n107), .Q(dataOut[21]) );
  DFFASRX1 \dataOut_reg[20]  ( .D(N273), .CLK(clk_out), .RSTB(n74), .SETB(n106), .Q(dataOut[20]) );
  DFFASRX1 \dataOut_reg[19]  ( .D(N272), .CLK(clk_out), .RSTB(n73), .SETB(n105), .Q(dataOut[19]) );
  DFFASRX1 \dataOut_reg[18]  ( .D(N271), .CLK(clk_out), .RSTB(n72), .SETB(n104), .Q(dataOut[18]) );
  DFFASRX1 \dataOut_reg[17]  ( .D(N270), .CLK(clk_out), .RSTB(n71), .SETB(n103), .Q(dataOut[17]) );
  DFFASRX1 \dataOut_reg[16]  ( .D(N269), .CLK(clk_out), .RSTB(n70), .SETB(n102), .Q(dataOut[16]) );
  DFFASRX1 \dataOut_reg[15]  ( .D(N268), .CLK(clk_out), .RSTB(n69), .SETB(n101), .Q(dataOut[15]) );
  DFFASRX1 \dataOut_reg[14]  ( .D(N267), .CLK(clk_out), .RSTB(n68), .SETB(n100), .Q(dataOut[14]) );
  DFFASRX1 \dataOut_reg[13]  ( .D(N266), .CLK(clk_out), .RSTB(n67), .SETB(n99), 
        .Q(dataOut[13]) );
  DFFASRX1 \dataOut_reg[12]  ( .D(N265), .CLK(clk_out), .RSTB(n66), .SETB(n98), 
        .Q(dataOut[12]) );
  DFFASRX1 \dataOut_reg[11]  ( .D(N264), .CLK(clk_out), .RSTB(n65), .SETB(n97), 
        .Q(dataOut[11]) );
  DFFASRX1 \dataOut_reg[10]  ( .D(N263), .CLK(clk_out), .RSTB(n64), .SETB(n96), 
        .Q(dataOut[10]) );
  DFFASRX1 \dataOut_reg[9]  ( .D(N262), .CLK(clk_out), .RSTB(n63), .SETB(n95), 
        .Q(dataOut[9]) );
  DFFASRX1 \dataOut_reg[8]  ( .D(N261), .CLK(clk_out), .RSTB(n62), .SETB(n94), 
        .Q(dataOut[8]) );
  DFFASRX1 \dataOut_reg[7]  ( .D(N260), .CLK(clk_out), .RSTB(n61), .SETB(n93), 
        .Q(dataOut[7]) );
  DFFASRX1 \dataOut_reg[6]  ( .D(N259), .CLK(clk_out), .RSTB(n60), .SETB(n92), 
        .Q(dataOut[6]) );
  DFFASRX1 \dataOut_reg[5]  ( .D(N258), .CLK(clk_out), .RSTB(n59), .SETB(n91), 
        .Q(dataOut[5]) );
  DFFASRX1 \dataOut_reg[4]  ( .D(N257), .CLK(clk_out), .RSTB(n58), .SETB(n90), 
        .Q(dataOut[4]) );
  DFFASRX1 \dataOut_reg[3]  ( .D(N256), .CLK(clk_out), .RSTB(n57), .SETB(n89), 
        .Q(dataOut[3]) );
  DFFASRX1 \dataOut_reg[2]  ( .D(N255), .CLK(clk_out), .RSTB(n56), .SETB(n88), 
        .Q(dataOut[2]) );
  DFFASRX1 \dataOut_reg[1]  ( .D(N254), .CLK(clk_out), .RSTB(n55), .SETB(n87), 
        .Q(dataOut[1]) );
  DFFASRX1 \dataOut_reg[0]  ( .D(N253), .CLK(clk_out), .RSTB(n54), .SETB(n86), 
        .Q(dataOut[0]) );
  AO22X1 U306 ( .IN1(n6828), .IN2(n7083), .IN3(\FIFO[127][24] ), .IN4(n7087), 
        .Q(n491) );
  AO22X1 U307 ( .IN1(n6817), .IN2(n7084), .IN3(\FIFO[127][25] ), .IN4(n7087), 
        .Q(n492) );
  AO22X1 U308 ( .IN1(n6806), .IN2(n206), .IN3(\FIFO[127][26] ), .IN4(n7087), 
        .Q(n493) );
  AO22X1 U309 ( .IN1(n6795), .IN2(n206), .IN3(\FIFO[127][27] ), .IN4(n7087), 
        .Q(n494) );
  AO22X1 U310 ( .IN1(n6784), .IN2(n7084), .IN3(\FIFO[127][28] ), .IN4(n7087), 
        .Q(n495) );
  AO22X1 U311 ( .IN1(n6773), .IN2(n7083), .IN3(\FIFO[127][29] ), .IN4(n7087), 
        .Q(n496) );
  AO22X1 U312 ( .IN1(n6762), .IN2(n7082), .IN3(\FIFO[127][30] ), .IN4(n7087), 
        .Q(n497) );
  AO22X1 U313 ( .IN1(n6751), .IN2(n206), .IN3(\FIFO[127][31] ), .IN4(n7087), 
        .Q(n498) );
  AO21X1 U314 ( .IN1(n238), .IN2(n239), .IN3(n5974), .Q(n206) );
  AO22X1 U339 ( .IN1(n6828), .IN2(n6737), .IN3(\FIFO[126][24] ), .IN4(n6740), 
        .Q(n523) );
  AO22X1 U340 ( .IN1(n6817), .IN2(n6735), .IN3(\FIFO[126][25] ), .IN4(n6740), 
        .Q(n524) );
  AO22X1 U341 ( .IN1(n6806), .IN2(n6736), .IN3(\FIFO[126][26] ), .IN4(n6740), 
        .Q(n525) );
  AO22X1 U342 ( .IN1(n6795), .IN2(n6737), .IN3(\FIFO[126][27] ), .IN4(n6740), 
        .Q(n526) );
  AO22X1 U343 ( .IN1(n6784), .IN2(n6736), .IN3(\FIFO[126][28] ), .IN4(n6740), 
        .Q(n527) );
  AO22X1 U344 ( .IN1(n6773), .IN2(n6735), .IN3(\FIFO[126][29] ), .IN4(n6740), 
        .Q(n528) );
  AO22X1 U345 ( .IN1(n6762), .IN2(n6737), .IN3(\FIFO[126][30] ), .IN4(n6740), 
        .Q(n529) );
  AO22X1 U346 ( .IN1(n6751), .IN2(n6736), .IN3(\FIFO[126][31] ), .IN4(n6740), 
        .Q(n530) );
  AO21X1 U347 ( .IN1(n241), .IN2(n239), .IN3(n5975), .Q(n240) );
  AO22X1 U372 ( .IN1(n6828), .IN2(n6729), .IN3(\FIFO[125][24] ), .IN4(n6734), 
        .Q(n555) );
  AO22X1 U373 ( .IN1(n6817), .IN2(n6729), .IN3(\FIFO[125][25] ), .IN4(n6734), 
        .Q(n556) );
  AO22X1 U374 ( .IN1(n6806), .IN2(n6729), .IN3(\FIFO[125][26] ), .IN4(n6734), 
        .Q(n557) );
  AO22X1 U375 ( .IN1(n6795), .IN2(n6729), .IN3(\FIFO[125][27] ), .IN4(n6734), 
        .Q(n558) );
  AO22X1 U376 ( .IN1(n6784), .IN2(n6730), .IN3(\FIFO[125][28] ), .IN4(n6734), 
        .Q(n559) );
  AO22X1 U377 ( .IN1(n6773), .IN2(n6729), .IN3(\FIFO[125][29] ), .IN4(n6734), 
        .Q(n560) );
  AO22X1 U378 ( .IN1(n6762), .IN2(n6731), .IN3(\FIFO[125][30] ), .IN4(n6734), 
        .Q(n561) );
  AO22X1 U379 ( .IN1(n6751), .IN2(n6730), .IN3(\FIFO[125][31] ), .IN4(n6734), 
        .Q(n562) );
  AO21X1 U380 ( .IN1(n243), .IN2(n239), .IN3(n5974), .Q(n242) );
  AO22X1 U393 ( .IN1(n6960), .IN2(n6724), .IN3(\FIFO[124][12] ), .IN4(n6727), 
        .Q(n575) );
  AO22X1 U394 ( .IN1(n6949), .IN2(n6724), .IN3(\FIFO[124][13] ), .IN4(n6727), 
        .Q(n576) );
  AO22X1 U395 ( .IN1(n6938), .IN2(n6723), .IN3(\FIFO[124][14] ), .IN4(n6727), 
        .Q(n577) );
  AO22X1 U396 ( .IN1(n6927), .IN2(n6723), .IN3(\FIFO[124][15] ), .IN4(n6727), 
        .Q(n578) );
  AO22X1 U397 ( .IN1(n6916), .IN2(n6723), .IN3(\FIFO[124][16] ), .IN4(n6727), 
        .Q(n579) );
  AO22X1 U398 ( .IN1(n6905), .IN2(n6723), .IN3(\FIFO[124][17] ), .IN4(n6727), 
        .Q(n580) );
  AO22X1 U405 ( .IN1(n6828), .IN2(n244), .IN3(\FIFO[124][24] ), .IN4(n6728), 
        .Q(n587) );
  AO22X1 U406 ( .IN1(n6817), .IN2(n244), .IN3(\FIFO[124][25] ), .IN4(n6728), 
        .Q(n588) );
  AO22X1 U407 ( .IN1(n6806), .IN2(n244), .IN3(\FIFO[124][26] ), .IN4(n6728), 
        .Q(n589) );
  AO22X1 U408 ( .IN1(n6795), .IN2(n6725), .IN3(\FIFO[124][27] ), .IN4(n6728), 
        .Q(n590) );
  AO22X1 U409 ( .IN1(n6784), .IN2(n6725), .IN3(\FIFO[124][28] ), .IN4(n6728), 
        .Q(n591) );
  AO22X1 U410 ( .IN1(n6773), .IN2(n6724), .IN3(\FIFO[124][29] ), .IN4(n6728), 
        .Q(n592) );
  AO22X1 U411 ( .IN1(n6762), .IN2(n6723), .IN3(\FIFO[124][30] ), .IN4(n6728), 
        .Q(n593) );
  AO22X1 U412 ( .IN1(n6751), .IN2(n6724), .IN3(\FIFO[124][31] ), .IN4(n6728), 
        .Q(n594) );
  AO21X1 U413 ( .IN1(n245), .IN2(n239), .IN3(n5975), .Q(n244) );
  AO22X1 U438 ( .IN1(n6828), .IN2(n246), .IN3(\FIFO[123][24] ), .IN4(n6722), 
        .Q(n619) );
  AO22X1 U439 ( .IN1(n6817), .IN2(n246), .IN3(\FIFO[123][25] ), .IN4(n6722), 
        .Q(n620) );
  AO22X1 U440 ( .IN1(n6806), .IN2(n6717), .IN3(\FIFO[123][26] ), .IN4(n6722), 
        .Q(n621) );
  AO22X1 U441 ( .IN1(n6795), .IN2(n6718), .IN3(\FIFO[123][27] ), .IN4(n6722), 
        .Q(n622) );
  AO22X1 U442 ( .IN1(n6784), .IN2(n6719), .IN3(\FIFO[123][28] ), .IN4(n6722), 
        .Q(n623) );
  AO22X1 U443 ( .IN1(n6773), .IN2(n6719), .IN3(\FIFO[123][29] ), .IN4(n6722), 
        .Q(n624) );
  AO22X1 U444 ( .IN1(n6762), .IN2(n6718), .IN3(\FIFO[123][30] ), .IN4(n6722), 
        .Q(n625) );
  AO22X1 U445 ( .IN1(n6751), .IN2(n6717), .IN3(\FIFO[123][31] ), .IN4(n6722), 
        .Q(n626) );
  AO21X1 U446 ( .IN1(n247), .IN2(n239), .IN3(n5974), .Q(n246) );
  AO22X1 U471 ( .IN1(n6828), .IN2(n6712), .IN3(\FIFO[122][24] ), .IN4(n6716), 
        .Q(n651) );
  AO22X1 U472 ( .IN1(n6817), .IN2(n6713), .IN3(\FIFO[122][25] ), .IN4(n6716), 
        .Q(n652) );
  AO22X1 U473 ( .IN1(n6806), .IN2(n248), .IN3(\FIFO[122][26] ), .IN4(n6716), 
        .Q(n653) );
  AO22X1 U474 ( .IN1(n6795), .IN2(n248), .IN3(\FIFO[122][27] ), .IN4(n6716), 
        .Q(n654) );
  AO22X1 U475 ( .IN1(n6784), .IN2(n6713), .IN3(\FIFO[122][28] ), .IN4(n6716), 
        .Q(n655) );
  AO22X1 U476 ( .IN1(n6773), .IN2(n6712), .IN3(\FIFO[122][29] ), .IN4(n6716), 
        .Q(n656) );
  AO22X1 U477 ( .IN1(n6762), .IN2(n6711), .IN3(\FIFO[122][30] ), .IN4(n6716), 
        .Q(n657) );
  AO22X1 U478 ( .IN1(n6751), .IN2(n248), .IN3(\FIFO[122][31] ), .IN4(n6716), 
        .Q(n658) );
  AO21X1 U479 ( .IN1(n249), .IN2(n239), .IN3(n5975), .Q(n248) );
  AO22X1 U480 ( .IN1(n7098), .IN2(n6707), .IN3(\FIFO[121][0] ), .IN4(n6708), 
        .Q(n659) );
  AO22X1 U481 ( .IN1(n7081), .IN2(n6707), .IN3(\FIFO[121][1] ), .IN4(n6708), 
        .Q(n660) );
  AO22X1 U482 ( .IN1(n7070), .IN2(n6707), .IN3(\FIFO[121][2] ), .IN4(n6708), 
        .Q(n661) );
  AO22X1 U483 ( .IN1(n7059), .IN2(n6707), .IN3(\FIFO[121][3] ), .IN4(n6708), 
        .Q(n662) );
  AO22X1 U484 ( .IN1(n7048), .IN2(n6707), .IN3(\FIFO[121][4] ), .IN4(n6708), 
        .Q(n663) );
  AO22X1 U485 ( .IN1(n7037), .IN2(n6707), .IN3(\FIFO[121][5] ), .IN4(n6708), 
        .Q(n664) );
  AO22X1 U486 ( .IN1(n7026), .IN2(n6707), .IN3(\FIFO[121][6] ), .IN4(n6708), 
        .Q(n665) );
  AO22X1 U487 ( .IN1(n7015), .IN2(n6706), .IN3(\FIFO[121][7] ), .IN4(n6708), 
        .Q(n666) );
  AO22X1 U488 ( .IN1(n7004), .IN2(n6706), .IN3(\FIFO[121][8] ), .IN4(n6708), 
        .Q(n667) );
  AO22X1 U489 ( .IN1(n6993), .IN2(n6706), .IN3(\FIFO[121][9] ), .IN4(n6708), 
        .Q(n668) );
  AO22X1 U490 ( .IN1(n6982), .IN2(n6706), .IN3(\FIFO[121][10] ), .IN4(n6708), 
        .Q(n669) );
  AO22X1 U491 ( .IN1(n6971), .IN2(n6706), .IN3(\FIFO[121][11] ), .IN4(n6708), 
        .Q(n670) );
  AO22X1 U492 ( .IN1(n6960), .IN2(n6706), .IN3(\FIFO[121][12] ), .IN4(n6709), 
        .Q(n671) );
  AO22X1 U493 ( .IN1(n6949), .IN2(n6706), .IN3(\FIFO[121][13] ), .IN4(n6709), 
        .Q(n672) );
  AO22X1 U494 ( .IN1(n6938), .IN2(n6705), .IN3(\FIFO[121][14] ), .IN4(n6709), 
        .Q(n673) );
  AO22X1 U495 ( .IN1(n6927), .IN2(n6705), .IN3(\FIFO[121][15] ), .IN4(n6709), 
        .Q(n674) );
  AO22X1 U496 ( .IN1(n6916), .IN2(n6705), .IN3(\FIFO[121][16] ), .IN4(n6709), 
        .Q(n675) );
  AO22X1 U497 ( .IN1(n6905), .IN2(n6705), .IN3(\FIFO[121][17] ), .IN4(n6709), 
        .Q(n676) );
  AO22X1 U498 ( .IN1(n6894), .IN2(n6705), .IN3(\FIFO[121][18] ), .IN4(n6709), 
        .Q(n677) );
  AO22X1 U499 ( .IN1(n6883), .IN2(n6705), .IN3(\FIFO[121][19] ), .IN4(n6709), 
        .Q(n678) );
  AO22X1 U500 ( .IN1(n6872), .IN2(n6705), .IN3(\FIFO[121][20] ), .IN4(n6709), 
        .Q(n679) );
  AO22X1 U501 ( .IN1(n6861), .IN2(n6707), .IN3(\FIFO[121][21] ), .IN4(n6709), 
        .Q(n680) );
  AO22X1 U502 ( .IN1(n6850), .IN2(n6706), .IN3(\FIFO[121][22] ), .IN4(n6709), 
        .Q(n681) );
  AO22X1 U503 ( .IN1(n6839), .IN2(n6705), .IN3(\FIFO[121][23] ), .IN4(n6709), 
        .Q(n682) );
  AO22X1 U504 ( .IN1(n6828), .IN2(n250), .IN3(\FIFO[121][24] ), .IN4(n6710), 
        .Q(n683) );
  AO22X1 U505 ( .IN1(n6817), .IN2(n250), .IN3(\FIFO[121][25] ), .IN4(n6710), 
        .Q(n684) );
  AO22X1 U506 ( .IN1(n6806), .IN2(n250), .IN3(\FIFO[121][26] ), .IN4(n6710), 
        .Q(n685) );
  AO22X1 U507 ( .IN1(n6795), .IN2(n6707), .IN3(\FIFO[121][27] ), .IN4(n6710), 
        .Q(n686) );
  AO22X1 U508 ( .IN1(n6784), .IN2(n6706), .IN3(\FIFO[121][28] ), .IN4(n6710), 
        .Q(n687) );
  AO22X1 U509 ( .IN1(n6773), .IN2(n6707), .IN3(\FIFO[121][29] ), .IN4(n6710), 
        .Q(n688) );
  AO22X1 U510 ( .IN1(n6762), .IN2(n6706), .IN3(\FIFO[121][30] ), .IN4(n6710), 
        .Q(n689) );
  AO22X1 U511 ( .IN1(n6751), .IN2(n6705), .IN3(\FIFO[121][31] ), .IN4(n6710), 
        .Q(n690) );
  AO21X1 U512 ( .IN1(n251), .IN2(n239), .IN3(n5974), .Q(n250) );
  AO22X1 U513 ( .IN1(n7098), .IN2(n6701), .IN3(\FIFO[120][0] ), .IN4(n6702), 
        .Q(n691) );
  AO22X1 U514 ( .IN1(n7081), .IN2(n6701), .IN3(\FIFO[120][1] ), .IN4(n6702), 
        .Q(n692) );
  AO22X1 U515 ( .IN1(n7070), .IN2(n6701), .IN3(\FIFO[120][2] ), .IN4(n6702), 
        .Q(n693) );
  AO22X1 U516 ( .IN1(n7059), .IN2(n6701), .IN3(\FIFO[120][3] ), .IN4(n6702), 
        .Q(n694) );
  AO22X1 U517 ( .IN1(n7048), .IN2(n6701), .IN3(\FIFO[120][4] ), .IN4(n6702), 
        .Q(n695) );
  AO22X1 U518 ( .IN1(n7037), .IN2(n6701), .IN3(\FIFO[120][5] ), .IN4(n6702), 
        .Q(n696) );
  AO22X1 U519 ( .IN1(n7026), .IN2(n6701), .IN3(\FIFO[120][6] ), .IN4(n6702), 
        .Q(n697) );
  AO22X1 U520 ( .IN1(n7015), .IN2(n6700), .IN3(\FIFO[120][7] ), .IN4(n6702), 
        .Q(n698) );
  AO22X1 U521 ( .IN1(n7004), .IN2(n6700), .IN3(\FIFO[120][8] ), .IN4(n6702), 
        .Q(n699) );
  AO22X1 U522 ( .IN1(n6993), .IN2(n6700), .IN3(\FIFO[120][9] ), .IN4(n6702), 
        .Q(n700) );
  AO22X1 U523 ( .IN1(n6982), .IN2(n6700), .IN3(\FIFO[120][10] ), .IN4(n6702), 
        .Q(n701) );
  AO22X1 U524 ( .IN1(n6971), .IN2(n6700), .IN3(\FIFO[120][11] ), .IN4(n6702), 
        .Q(n702) );
  AO22X1 U525 ( .IN1(n6960), .IN2(n6700), .IN3(\FIFO[120][12] ), .IN4(n6703), 
        .Q(n703) );
  AO22X1 U526 ( .IN1(n6949), .IN2(n6700), .IN3(\FIFO[120][13] ), .IN4(n6703), 
        .Q(n704) );
  AO22X1 U527 ( .IN1(n6938), .IN2(n6699), .IN3(\FIFO[120][14] ), .IN4(n6703), 
        .Q(n705) );
  AO22X1 U528 ( .IN1(n6927), .IN2(n6699), .IN3(\FIFO[120][15] ), .IN4(n6703), 
        .Q(n706) );
  AO22X1 U529 ( .IN1(n6916), .IN2(n6699), .IN3(\FIFO[120][16] ), .IN4(n6703), 
        .Q(n707) );
  AO22X1 U530 ( .IN1(n6905), .IN2(n6699), .IN3(\FIFO[120][17] ), .IN4(n6703), 
        .Q(n708) );
  AO22X1 U531 ( .IN1(n6894), .IN2(n6699), .IN3(\FIFO[120][18] ), .IN4(n6703), 
        .Q(n709) );
  AO22X1 U532 ( .IN1(n6883), .IN2(n6699), .IN3(\FIFO[120][19] ), .IN4(n6703), 
        .Q(n710) );
  AO22X1 U533 ( .IN1(n6872), .IN2(n6699), .IN3(\FIFO[120][20] ), .IN4(n6703), 
        .Q(n711) );
  AO22X1 U534 ( .IN1(n6861), .IN2(n6701), .IN3(\FIFO[120][21] ), .IN4(n6703), 
        .Q(n712) );
  AO22X1 U535 ( .IN1(n6850), .IN2(n6700), .IN3(\FIFO[120][22] ), .IN4(n6703), 
        .Q(n713) );
  AO22X1 U536 ( .IN1(n6839), .IN2(n6699), .IN3(\FIFO[120][23] ), .IN4(n6703), 
        .Q(n714) );
  AO22X1 U537 ( .IN1(n6828), .IN2(n252), .IN3(\FIFO[120][24] ), .IN4(n6704), 
        .Q(n715) );
  AO22X1 U538 ( .IN1(n6817), .IN2(n252), .IN3(\FIFO[120][25] ), .IN4(n6704), 
        .Q(n716) );
  AO22X1 U539 ( .IN1(n6806), .IN2(n252), .IN3(\FIFO[120][26] ), .IN4(n6704), 
        .Q(n717) );
  AO22X1 U540 ( .IN1(n6795), .IN2(n6701), .IN3(\FIFO[120][27] ), .IN4(n6704), 
        .Q(n718) );
  AO22X1 U541 ( .IN1(n6784), .IN2(n6700), .IN3(\FIFO[120][28] ), .IN4(n6704), 
        .Q(n719) );
  AO22X1 U542 ( .IN1(n6773), .IN2(n6701), .IN3(\FIFO[120][29] ), .IN4(n6704), 
        .Q(n720) );
  AO22X1 U543 ( .IN1(n6762), .IN2(n6700), .IN3(\FIFO[120][30] ), .IN4(n6704), 
        .Q(n721) );
  AO22X1 U544 ( .IN1(n6751), .IN2(n6699), .IN3(\FIFO[120][31] ), .IN4(n6704), 
        .Q(n722) );
  AO21X1 U545 ( .IN1(n253), .IN2(n239), .IN3(n5975), .Q(n252) );
  AO22X1 U570 ( .IN1(n6827), .IN2(n6693), .IN3(\FIFO[119][24] ), .IN4(n6698), 
        .Q(n747) );
  AO22X1 U571 ( .IN1(n6816), .IN2(n6693), .IN3(\FIFO[119][25] ), .IN4(n6698), 
        .Q(n748) );
  AO22X1 U572 ( .IN1(n6805), .IN2(n6693), .IN3(\FIFO[119][26] ), .IN4(n6698), 
        .Q(n749) );
  AO22X1 U573 ( .IN1(n6794), .IN2(n6693), .IN3(\FIFO[119][27] ), .IN4(n6698), 
        .Q(n750) );
  AO22X1 U574 ( .IN1(n6783), .IN2(n6693), .IN3(\FIFO[119][28] ), .IN4(n6698), 
        .Q(n751) );
  AO22X1 U575 ( .IN1(n6772), .IN2(n6694), .IN3(\FIFO[119][29] ), .IN4(n6698), 
        .Q(n752) );
  AO22X1 U576 ( .IN1(n6761), .IN2(n6693), .IN3(\FIFO[119][30] ), .IN4(n6698), 
        .Q(n753) );
  AO22X1 U577 ( .IN1(n6750), .IN2(n6694), .IN3(\FIFO[119][31] ), .IN4(n6698), 
        .Q(n754) );
  AO21X1 U578 ( .IN1(n255), .IN2(n239), .IN3(n5974), .Q(n254) );
  AO22X1 U603 ( .IN1(n6827), .IN2(n256), .IN3(\FIFO[118][24] ), .IN4(n6692), 
        .Q(n779) );
  AO22X1 U604 ( .IN1(n6816), .IN2(n256), .IN3(\FIFO[118][25] ), .IN4(n6692), 
        .Q(n780) );
  AO22X1 U605 ( .IN1(n6805), .IN2(n6687), .IN3(\FIFO[118][26] ), .IN4(n6692), 
        .Q(n781) );
  AO22X1 U606 ( .IN1(n6794), .IN2(n6688), .IN3(\FIFO[118][27] ), .IN4(n6692), 
        .Q(n782) );
  AO22X1 U607 ( .IN1(n6783), .IN2(n6689), .IN3(\FIFO[118][28] ), .IN4(n6692), 
        .Q(n783) );
  AO22X1 U608 ( .IN1(n6772), .IN2(n6689), .IN3(\FIFO[118][29] ), .IN4(n6692), 
        .Q(n784) );
  AO22X1 U609 ( .IN1(n6761), .IN2(n6688), .IN3(\FIFO[118][30] ), .IN4(n6692), 
        .Q(n785) );
  AO22X1 U610 ( .IN1(n6750), .IN2(n6687), .IN3(\FIFO[118][31] ), .IN4(n6692), 
        .Q(n786) );
  AO21X1 U611 ( .IN1(n257), .IN2(n239), .IN3(n5975), .Q(n256) );
  AO22X1 U612 ( .IN1(n7097), .IN2(n6683), .IN3(\FIFO[117][0] ), .IN4(n6684), 
        .Q(n787) );
  AO22X1 U613 ( .IN1(n7080), .IN2(n6682), .IN3(\FIFO[117][1] ), .IN4(n6684), 
        .Q(n788) );
  AO22X1 U614 ( .IN1(n7069), .IN2(n6681), .IN3(\FIFO[117][2] ), .IN4(n6684), 
        .Q(n789) );
  AO22X1 U615 ( .IN1(n7058), .IN2(n6683), .IN3(\FIFO[117][3] ), .IN4(n6684), 
        .Q(n790) );
  AO22X1 U616 ( .IN1(n7047), .IN2(n6682), .IN3(\FIFO[117][4] ), .IN4(n6684), 
        .Q(n791) );
  AO22X1 U617 ( .IN1(n7036), .IN2(n6681), .IN3(\FIFO[117][5] ), .IN4(n6684), 
        .Q(n792) );
  AO22X1 U618 ( .IN1(n7025), .IN2(n6683), .IN3(\FIFO[117][6] ), .IN4(n6684), 
        .Q(n793) );
  AO22X1 U619 ( .IN1(n7014), .IN2(n6683), .IN3(\FIFO[117][7] ), .IN4(n6684), 
        .Q(n794) );
  AO22X1 U620 ( .IN1(n7003), .IN2(n6683), .IN3(\FIFO[117][8] ), .IN4(n6684), 
        .Q(n795) );
  AO22X1 U621 ( .IN1(n6992), .IN2(n6683), .IN3(\FIFO[117][9] ), .IN4(n6684), 
        .Q(n796) );
  AO22X1 U622 ( .IN1(n6981), .IN2(n6683), .IN3(\FIFO[117][10] ), .IN4(n6684), 
        .Q(n797) );
  AO22X1 U623 ( .IN1(n6970), .IN2(n6683), .IN3(\FIFO[117][11] ), .IN4(n6684), 
        .Q(n798) );
  AO22X1 U624 ( .IN1(n6959), .IN2(n6683), .IN3(\FIFO[117][12] ), .IN4(n6685), 
        .Q(n799) );
  AO22X1 U625 ( .IN1(n6948), .IN2(n6683), .IN3(\FIFO[117][13] ), .IN4(n6685), 
        .Q(n800) );
  AO22X1 U626 ( .IN1(n6937), .IN2(n6682), .IN3(\FIFO[117][14] ), .IN4(n6685), 
        .Q(n801) );
  AO22X1 U627 ( .IN1(n6926), .IN2(n6682), .IN3(\FIFO[117][15] ), .IN4(n6685), 
        .Q(n802) );
  AO22X1 U628 ( .IN1(n6915), .IN2(n6682), .IN3(\FIFO[117][16] ), .IN4(n6685), 
        .Q(n803) );
  AO22X1 U629 ( .IN1(n6904), .IN2(n6682), .IN3(\FIFO[117][17] ), .IN4(n6685), 
        .Q(n804) );
  AO22X1 U630 ( .IN1(n6893), .IN2(n6682), .IN3(\FIFO[117][18] ), .IN4(n6685), 
        .Q(n805) );
  AO22X1 U631 ( .IN1(n6882), .IN2(n6682), .IN3(\FIFO[117][19] ), .IN4(n6685), 
        .Q(n806) );
  AO22X1 U632 ( .IN1(n6871), .IN2(n6682), .IN3(\FIFO[117][20] ), .IN4(n6685), 
        .Q(n807) );
  AO22X1 U633 ( .IN1(n6860), .IN2(n6681), .IN3(\FIFO[117][21] ), .IN4(n6685), 
        .Q(n808) );
  AO22X1 U634 ( .IN1(n6849), .IN2(n6681), .IN3(\FIFO[117][22] ), .IN4(n6685), 
        .Q(n809) );
  AO22X1 U635 ( .IN1(n6838), .IN2(n6681), .IN3(\FIFO[117][23] ), .IN4(n6685), 
        .Q(n810) );
  AO22X1 U636 ( .IN1(n6827), .IN2(n6681), .IN3(\FIFO[117][24] ), .IN4(n6686), 
        .Q(n811) );
  AO22X1 U637 ( .IN1(n6816), .IN2(n6681), .IN3(\FIFO[117][25] ), .IN4(n6686), 
        .Q(n812) );
  AO22X1 U638 ( .IN1(n6805), .IN2(n6681), .IN3(\FIFO[117][26] ), .IN4(n6686), 
        .Q(n813) );
  AO22X1 U639 ( .IN1(n6794), .IN2(n6681), .IN3(\FIFO[117][27] ), .IN4(n6686), 
        .Q(n814) );
  AO22X1 U640 ( .IN1(n6783), .IN2(n6681), .IN3(\FIFO[117][28] ), .IN4(n6686), 
        .Q(n815) );
  AO22X1 U641 ( .IN1(n6772), .IN2(n6682), .IN3(\FIFO[117][29] ), .IN4(n6686), 
        .Q(n816) );
  AO22X1 U642 ( .IN1(n6761), .IN2(n6681), .IN3(\FIFO[117][30] ), .IN4(n6686), 
        .Q(n817) );
  AO22X1 U643 ( .IN1(n6750), .IN2(n6682), .IN3(\FIFO[117][31] ), .IN4(n6686), 
        .Q(n818) );
  AO21X1 U644 ( .IN1(n259), .IN2(n239), .IN3(n5974), .Q(n258) );
  AO22X1 U645 ( .IN1(n7097), .IN2(n6677), .IN3(\FIFO[116][0] ), .IN4(n6678), 
        .Q(n819) );
  AO22X1 U646 ( .IN1(n7080), .IN2(n6677), .IN3(\FIFO[116][1] ), .IN4(n6678), 
        .Q(n820) );
  AO22X1 U647 ( .IN1(n7069), .IN2(n6677), .IN3(\FIFO[116][2] ), .IN4(n6678), 
        .Q(n821) );
  AO22X1 U648 ( .IN1(n7058), .IN2(n6677), .IN3(\FIFO[116][3] ), .IN4(n6678), 
        .Q(n822) );
  AO22X1 U649 ( .IN1(n7047), .IN2(n6677), .IN3(\FIFO[116][4] ), .IN4(n6678), 
        .Q(n823) );
  AO22X1 U650 ( .IN1(n7036), .IN2(n6677), .IN3(\FIFO[116][5] ), .IN4(n6678), 
        .Q(n824) );
  AO22X1 U651 ( .IN1(n7025), .IN2(n6677), .IN3(\FIFO[116][6] ), .IN4(n6678), 
        .Q(n825) );
  AO22X1 U652 ( .IN1(n7014), .IN2(n6676), .IN3(\FIFO[116][7] ), .IN4(n6678), 
        .Q(n826) );
  AO22X1 U653 ( .IN1(n7003), .IN2(n6676), .IN3(\FIFO[116][8] ), .IN4(n6678), 
        .Q(n827) );
  AO22X1 U654 ( .IN1(n6992), .IN2(n6676), .IN3(\FIFO[116][9] ), .IN4(n6678), 
        .Q(n828) );
  AO22X1 U655 ( .IN1(n6981), .IN2(n6676), .IN3(\FIFO[116][10] ), .IN4(n6678), 
        .Q(n829) );
  AO22X1 U656 ( .IN1(n6970), .IN2(n6676), .IN3(\FIFO[116][11] ), .IN4(n6678), 
        .Q(n830) );
  AO22X1 U657 ( .IN1(n6959), .IN2(n6676), .IN3(\FIFO[116][12] ), .IN4(n6679), 
        .Q(n831) );
  AO22X1 U658 ( .IN1(n6948), .IN2(n6676), .IN3(\FIFO[116][13] ), .IN4(n6679), 
        .Q(n832) );
  AO22X1 U659 ( .IN1(n6937), .IN2(n6675), .IN3(\FIFO[116][14] ), .IN4(n6679), 
        .Q(n833) );
  AO22X1 U660 ( .IN1(n6926), .IN2(n6675), .IN3(\FIFO[116][15] ), .IN4(n6679), 
        .Q(n834) );
  AO22X1 U661 ( .IN1(n6915), .IN2(n6675), .IN3(\FIFO[116][16] ), .IN4(n6679), 
        .Q(n835) );
  AO22X1 U662 ( .IN1(n6904), .IN2(n6675), .IN3(\FIFO[116][17] ), .IN4(n6679), 
        .Q(n836) );
  AO22X1 U663 ( .IN1(n6893), .IN2(n6675), .IN3(\FIFO[116][18] ), .IN4(n6679), 
        .Q(n837) );
  AO22X1 U664 ( .IN1(n6882), .IN2(n6675), .IN3(\FIFO[116][19] ), .IN4(n6679), 
        .Q(n838) );
  AO22X1 U665 ( .IN1(n6871), .IN2(n6675), .IN3(\FIFO[116][20] ), .IN4(n6679), 
        .Q(n839) );
  AO22X1 U666 ( .IN1(n6860), .IN2(n6677), .IN3(\FIFO[116][21] ), .IN4(n6679), 
        .Q(n840) );
  AO22X1 U667 ( .IN1(n6849), .IN2(n6676), .IN3(\FIFO[116][22] ), .IN4(n6679), 
        .Q(n841) );
  AO22X1 U668 ( .IN1(n6838), .IN2(n6675), .IN3(\FIFO[116][23] ), .IN4(n6679), 
        .Q(n842) );
  AO22X1 U669 ( .IN1(n6827), .IN2(n260), .IN3(\FIFO[116][24] ), .IN4(n6680), 
        .Q(n843) );
  AO22X1 U670 ( .IN1(n6816), .IN2(n260), .IN3(\FIFO[116][25] ), .IN4(n6680), 
        .Q(n844) );
  AO22X1 U671 ( .IN1(n6805), .IN2(n260), .IN3(\FIFO[116][26] ), .IN4(n6680), 
        .Q(n845) );
  AO22X1 U672 ( .IN1(n6794), .IN2(n6677), .IN3(\FIFO[116][27] ), .IN4(n6680), 
        .Q(n846) );
  AO22X1 U673 ( .IN1(n6783), .IN2(n6676), .IN3(\FIFO[116][28] ), .IN4(n6680), 
        .Q(n847) );
  AO22X1 U674 ( .IN1(n6772), .IN2(n6677), .IN3(\FIFO[116][29] ), .IN4(n6680), 
        .Q(n848) );
  AO22X1 U675 ( .IN1(n6761), .IN2(n6676), .IN3(\FIFO[116][30] ), .IN4(n6680), 
        .Q(n849) );
  AO22X1 U676 ( .IN1(n6750), .IN2(n6675), .IN3(\FIFO[116][31] ), .IN4(n6680), 
        .Q(n850) );
  AO21X1 U677 ( .IN1(n261), .IN2(n239), .IN3(n5975), .Q(n260) );
  AO22X1 U702 ( .IN1(n6827), .IN2(n6669), .IN3(\FIFO[115][24] ), .IN4(n6674), 
        .Q(n875) );
  AO22X1 U703 ( .IN1(n6816), .IN2(n6669), .IN3(\FIFO[115][25] ), .IN4(n6674), 
        .Q(n876) );
  AO22X1 U704 ( .IN1(n6805), .IN2(n6669), .IN3(\FIFO[115][26] ), .IN4(n6674), 
        .Q(n877) );
  AO22X1 U705 ( .IN1(n6794), .IN2(n6669), .IN3(\FIFO[115][27] ), .IN4(n6674), 
        .Q(n878) );
  AO22X1 U706 ( .IN1(n6783), .IN2(n6670), .IN3(\FIFO[115][28] ), .IN4(n6674), 
        .Q(n879) );
  AO22X1 U707 ( .IN1(n6772), .IN2(n6669), .IN3(\FIFO[115][29] ), .IN4(n6674), 
        .Q(n880) );
  AO22X1 U708 ( .IN1(n6761), .IN2(n6671), .IN3(\FIFO[115][30] ), .IN4(n6674), 
        .Q(n881) );
  AO22X1 U709 ( .IN1(n6750), .IN2(n6670), .IN3(\FIFO[115][31] ), .IN4(n6674), 
        .Q(n882) );
  AO21X1 U710 ( .IN1(n263), .IN2(n239), .IN3(n5974), .Q(n262) );
  AO22X1 U735 ( .IN1(n6827), .IN2(n6663), .IN3(\FIFO[114][24] ), .IN4(n6668), 
        .Q(n907) );
  AO22X1 U736 ( .IN1(n6816), .IN2(n6663), .IN3(\FIFO[114][25] ), .IN4(n6668), 
        .Q(n908) );
  AO22X1 U737 ( .IN1(n6805), .IN2(n6663), .IN3(\FIFO[114][26] ), .IN4(n6668), 
        .Q(n909) );
  AO22X1 U738 ( .IN1(n6794), .IN2(n6663), .IN3(\FIFO[114][27] ), .IN4(n6668), 
        .Q(n910) );
  AO22X1 U739 ( .IN1(n6783), .IN2(n6663), .IN3(\FIFO[114][28] ), .IN4(n6668), 
        .Q(n911) );
  AO22X1 U740 ( .IN1(n6772), .IN2(n6664), .IN3(\FIFO[114][29] ), .IN4(n6668), 
        .Q(n912) );
  AO22X1 U741 ( .IN1(n6761), .IN2(n6663), .IN3(\FIFO[114][30] ), .IN4(n6668), 
        .Q(n913) );
  AO22X1 U742 ( .IN1(n6750), .IN2(n6664), .IN3(\FIFO[114][31] ), .IN4(n6668), 
        .Q(n914) );
  AO21X1 U743 ( .IN1(n265), .IN2(n239), .IN3(n5975), .Q(n264) );
  AO22X1 U744 ( .IN1(n7097), .IN2(n6659), .IN3(\FIFO[113][0] ), .IN4(n6660), 
        .Q(n915) );
  AO22X1 U745 ( .IN1(n7080), .IN2(n6659), .IN3(\FIFO[113][1] ), .IN4(n6660), 
        .Q(n916) );
  AO22X1 U746 ( .IN1(n7069), .IN2(n6659), .IN3(\FIFO[113][2] ), .IN4(n6660), 
        .Q(n917) );
  AO22X1 U747 ( .IN1(n7058), .IN2(n6659), .IN3(\FIFO[113][3] ), .IN4(n6660), 
        .Q(n918) );
  AO22X1 U748 ( .IN1(n7047), .IN2(n6659), .IN3(\FIFO[113][4] ), .IN4(n6660), 
        .Q(n919) );
  AO22X1 U749 ( .IN1(n7036), .IN2(n6659), .IN3(\FIFO[113][5] ), .IN4(n6660), 
        .Q(n920) );
  AO22X1 U750 ( .IN1(n7025), .IN2(n6659), .IN3(\FIFO[113][6] ), .IN4(n6660), 
        .Q(n921) );
  AO22X1 U752 ( .IN1(n7003), .IN2(n6658), .IN3(\FIFO[113][8] ), .IN4(n6660), 
        .Q(n923) );
  AO22X1 U753 ( .IN1(n6992), .IN2(n6658), .IN3(\FIFO[113][9] ), .IN4(n6660), 
        .Q(n924) );
  AO22X1 U754 ( .IN1(n6981), .IN2(n6658), .IN3(\FIFO[113][10] ), .IN4(n6660), 
        .Q(n925) );
  AO22X1 U755 ( .IN1(n6970), .IN2(n6658), .IN3(\FIFO[113][11] ), .IN4(n6660), 
        .Q(n926) );
  AO22X1 U756 ( .IN1(n6959), .IN2(n6658), .IN3(\FIFO[113][12] ), .IN4(n6661), 
        .Q(n927) );
  AO22X1 U757 ( .IN1(n6948), .IN2(n6658), .IN3(\FIFO[113][13] ), .IN4(n6661), 
        .Q(n928) );
  AO22X1 U758 ( .IN1(n6937), .IN2(n6659), .IN3(\FIFO[113][14] ), .IN4(n6661), 
        .Q(n929) );
  AO22X1 U759 ( .IN1(n6926), .IN2(n6658), .IN3(\FIFO[113][15] ), .IN4(n6661), 
        .Q(n930) );
  AO22X1 U760 ( .IN1(n6915), .IN2(n6657), .IN3(\FIFO[113][16] ), .IN4(n6661), 
        .Q(n931) );
  AO22X1 U761 ( .IN1(n6904), .IN2(n6659), .IN3(\FIFO[113][17] ), .IN4(n6661), 
        .Q(n932) );
  AO22X1 U762 ( .IN1(n6893), .IN2(n6658), .IN3(\FIFO[113][18] ), .IN4(n6661), 
        .Q(n933) );
  AO22X1 U763 ( .IN1(n6882), .IN2(n6657), .IN3(\FIFO[113][19] ), .IN4(n6661), 
        .Q(n934) );
  AO22X1 U764 ( .IN1(n6871), .IN2(n6659), .IN3(\FIFO[113][20] ), .IN4(n6661), 
        .Q(n935) );
  AO22X1 U765 ( .IN1(n6860), .IN2(n6657), .IN3(\FIFO[113][21] ), .IN4(n6661), 
        .Q(n936) );
  AO22X1 U766 ( .IN1(n6849), .IN2(n6657), .IN3(\FIFO[113][22] ), .IN4(n6661), 
        .Q(n937) );
  AO22X1 U767 ( .IN1(n6838), .IN2(n6657), .IN3(\FIFO[113][23] ), .IN4(n6661), 
        .Q(n938) );
  AO22X1 U768 ( .IN1(n6827), .IN2(n6657), .IN3(\FIFO[113][24] ), .IN4(n6662), 
        .Q(n939) );
  AO22X1 U769 ( .IN1(n6816), .IN2(n6657), .IN3(\FIFO[113][25] ), .IN4(n6662), 
        .Q(n940) );
  AO22X1 U770 ( .IN1(n6805), .IN2(n6657), .IN3(\FIFO[113][26] ), .IN4(n6662), 
        .Q(n941) );
  AO22X1 U771 ( .IN1(n6794), .IN2(n6657), .IN3(\FIFO[113][27] ), .IN4(n6662), 
        .Q(n942) );
  AO22X1 U772 ( .IN1(n6783), .IN2(n6657), .IN3(\FIFO[113][28] ), .IN4(n6662), 
        .Q(n943) );
  AO22X1 U773 ( .IN1(n6772), .IN2(n6658), .IN3(\FIFO[113][29] ), .IN4(n6662), 
        .Q(n944) );
  AO22X1 U774 ( .IN1(n6761), .IN2(n6657), .IN3(\FIFO[113][30] ), .IN4(n6662), 
        .Q(n945) );
  AO22X1 U775 ( .IN1(n6750), .IN2(n6658), .IN3(\FIFO[113][31] ), .IN4(n6662), 
        .Q(n946) );
  AO21X1 U776 ( .IN1(n267), .IN2(n239), .IN3(n5974), .Q(n266) );
  AO22X1 U777 ( .IN1(n7097), .IN2(n6653), .IN3(\FIFO[112][0] ), .IN4(n6654), 
        .Q(n947) );
  AO22X1 U778 ( .IN1(n7080), .IN2(n6652), .IN3(\FIFO[112][1] ), .IN4(n6654), 
        .Q(n948) );
  AO22X1 U779 ( .IN1(n7069), .IN2(n6651), .IN3(\FIFO[112][2] ), .IN4(n6654), 
        .Q(n949) );
  AO22X1 U780 ( .IN1(n7058), .IN2(n6653), .IN3(\FIFO[112][3] ), .IN4(n6654), 
        .Q(n950) );
  AO22X1 U781 ( .IN1(n7047), .IN2(n6652), .IN3(\FIFO[112][4] ), .IN4(n6654), 
        .Q(n951) );
  AO22X1 U782 ( .IN1(n7036), .IN2(n6651), .IN3(\FIFO[112][5] ), .IN4(n6654), 
        .Q(n952) );
  AO22X1 U783 ( .IN1(n7025), .IN2(n6653), .IN3(\FIFO[112][6] ), .IN4(n6654), 
        .Q(n953) );
  AO22X1 U784 ( .IN1(n7014), .IN2(n6653), .IN3(\FIFO[112][7] ), .IN4(n6654), 
        .Q(n954) );
  AO22X1 U785 ( .IN1(n7003), .IN2(n6653), .IN3(\FIFO[112][8] ), .IN4(n6654), 
        .Q(n955) );
  AO22X1 U786 ( .IN1(n6992), .IN2(n6653), .IN3(\FIFO[112][9] ), .IN4(n6654), 
        .Q(n956) );
  AO22X1 U787 ( .IN1(n6981), .IN2(n6653), .IN3(\FIFO[112][10] ), .IN4(n6654), 
        .Q(n957) );
  AO22X1 U788 ( .IN1(n6970), .IN2(n6653), .IN3(\FIFO[112][11] ), .IN4(n6654), 
        .Q(n958) );
  AO22X1 U789 ( .IN1(n6959), .IN2(n6653), .IN3(\FIFO[112][12] ), .IN4(n6655), 
        .Q(n959) );
  AO22X1 U790 ( .IN1(n6948), .IN2(n6653), .IN3(\FIFO[112][13] ), .IN4(n6655), 
        .Q(n960) );
  AO22X1 U791 ( .IN1(n6937), .IN2(n6652), .IN3(\FIFO[112][14] ), .IN4(n6655), 
        .Q(n961) );
  AO22X1 U792 ( .IN1(n6926), .IN2(n6652), .IN3(\FIFO[112][15] ), .IN4(n6655), 
        .Q(n962) );
  AO22X1 U793 ( .IN1(n6915), .IN2(n6652), .IN3(\FIFO[112][16] ), .IN4(n6655), 
        .Q(n963) );
  AO22X1 U794 ( .IN1(n6904), .IN2(n6652), .IN3(\FIFO[112][17] ), .IN4(n6655), 
        .Q(n964) );
  AO22X1 U795 ( .IN1(n6893), .IN2(n6652), .IN3(\FIFO[112][18] ), .IN4(n6655), 
        .Q(n965) );
  AO22X1 U796 ( .IN1(n6882), .IN2(n6652), .IN3(\FIFO[112][19] ), .IN4(n6655), 
        .Q(n966) );
  AO22X1 U797 ( .IN1(n6871), .IN2(n6652), .IN3(\FIFO[112][20] ), .IN4(n6655), 
        .Q(n967) );
  AO22X1 U798 ( .IN1(n6860), .IN2(n6651), .IN3(\FIFO[112][21] ), .IN4(n6655), 
        .Q(n968) );
  AO22X1 U799 ( .IN1(n6849), .IN2(n6651), .IN3(\FIFO[112][22] ), .IN4(n6655), 
        .Q(n969) );
  AO22X1 U800 ( .IN1(n6838), .IN2(n6651), .IN3(\FIFO[112][23] ), .IN4(n6655), 
        .Q(n970) );
  AO22X1 U801 ( .IN1(n6827), .IN2(n6651), .IN3(\FIFO[112][24] ), .IN4(n6656), 
        .Q(n971) );
  AO22X1 U802 ( .IN1(n6816), .IN2(n6651), .IN3(\FIFO[112][25] ), .IN4(n6656), 
        .Q(n972) );
  AO22X1 U803 ( .IN1(n6805), .IN2(n6651), .IN3(\FIFO[112][26] ), .IN4(n6656), 
        .Q(n973) );
  AO22X1 U804 ( .IN1(n6794), .IN2(n6651), .IN3(\FIFO[112][27] ), .IN4(n6656), 
        .Q(n974) );
  AO22X1 U805 ( .IN1(n6783), .IN2(n6651), .IN3(\FIFO[112][28] ), .IN4(n6656), 
        .Q(n975) );
  AO22X1 U806 ( .IN1(n6772), .IN2(n6652), .IN3(\FIFO[112][29] ), .IN4(n6656), 
        .Q(n976) );
  AO22X1 U807 ( .IN1(n6761), .IN2(n6651), .IN3(\FIFO[112][30] ), .IN4(n6656), 
        .Q(n977) );
  AO22X1 U808 ( .IN1(n6750), .IN2(n6652), .IN3(\FIFO[112][31] ), .IN4(n6656), 
        .Q(n978) );
  AO21X1 U809 ( .IN1(n269), .IN2(n239), .IN3(n5975), .Q(n268) );
  AO22X1 U835 ( .IN1(n6827), .IN2(n271), .IN3(\FIFO[111][24] ), .IN4(n6650), 
        .Q(n1003) );
  AO22X1 U836 ( .IN1(n6816), .IN2(n271), .IN3(\FIFO[111][25] ), .IN4(n6650), 
        .Q(n1004) );
  AO22X1 U837 ( .IN1(n6805), .IN2(n271), .IN3(\FIFO[111][26] ), .IN4(n6650), 
        .Q(n1005) );
  AO22X1 U838 ( .IN1(n6794), .IN2(n6647), .IN3(\FIFO[111][27] ), .IN4(n6650), 
        .Q(n1006) );
  AO22X1 U839 ( .IN1(n6783), .IN2(n6646), .IN3(\FIFO[111][28] ), .IN4(n6650), 
        .Q(n1007) );
  AO22X1 U840 ( .IN1(n6772), .IN2(n6647), .IN3(\FIFO[111][29] ), .IN4(n6650), 
        .Q(n1008) );
  AO22X1 U841 ( .IN1(n6761), .IN2(n6646), .IN3(\FIFO[111][30] ), .IN4(n6650), 
        .Q(n1009) );
  AO22X1 U842 ( .IN1(n6750), .IN2(n6645), .IN3(\FIFO[111][31] ), .IN4(n6650), 
        .Q(n1010) );
  AO21X1 U843 ( .IN1(n272), .IN2(n238), .IN3(n5974), .Q(n271) );
  AO22X1 U868 ( .IN1(n6827), .IN2(n273), .IN3(\FIFO[110][24] ), .IN4(n6644), 
        .Q(n1035) );
  AO22X1 U869 ( .IN1(n6816), .IN2(n273), .IN3(\FIFO[110][25] ), .IN4(n6644), 
        .Q(n1036) );
  AO22X1 U870 ( .IN1(n6805), .IN2(n273), .IN3(\FIFO[110][26] ), .IN4(n6644), 
        .Q(n1037) );
  AO22X1 U871 ( .IN1(n6794), .IN2(n6641), .IN3(\FIFO[110][27] ), .IN4(n6644), 
        .Q(n1038) );
  AO22X1 U872 ( .IN1(n6783), .IN2(n6640), .IN3(\FIFO[110][28] ), .IN4(n6644), 
        .Q(n1039) );
  AO22X1 U873 ( .IN1(n6772), .IN2(n6641), .IN3(\FIFO[110][29] ), .IN4(n6644), 
        .Q(n1040) );
  AO22X1 U874 ( .IN1(n6761), .IN2(n6640), .IN3(\FIFO[110][30] ), .IN4(n6644), 
        .Q(n1041) );
  AO22X1 U875 ( .IN1(n6750), .IN2(n6639), .IN3(\FIFO[110][31] ), .IN4(n6644), 
        .Q(n1042) );
  AO21X1 U876 ( .IN1(n272), .IN2(n241), .IN3(n5975), .Q(n273) );
  AO22X1 U877 ( .IN1(n7097), .IN2(n6635), .IN3(\FIFO[109][0] ), .IN4(n6636), 
        .Q(n1043) );
  AO22X1 U878 ( .IN1(n7080), .IN2(n6635), .IN3(\FIFO[109][1] ), .IN4(n6636), 
        .Q(n1044) );
  AO22X1 U879 ( .IN1(n7069), .IN2(n6635), .IN3(\FIFO[109][2] ), .IN4(n6636), 
        .Q(n1045) );
  AO22X1 U880 ( .IN1(n7058), .IN2(n6635), .IN3(\FIFO[109][3] ), .IN4(n6636), 
        .Q(n1046) );
  AO22X1 U881 ( .IN1(n7047), .IN2(n6635), .IN3(\FIFO[109][4] ), .IN4(n6636), 
        .Q(n1047) );
  AO22X1 U882 ( .IN1(n7036), .IN2(n6635), .IN3(\FIFO[109][5] ), .IN4(n6636), 
        .Q(n1048) );
  AO22X1 U883 ( .IN1(n7025), .IN2(n6635), .IN3(\FIFO[109][6] ), .IN4(n6636), 
        .Q(n1049) );
  AO22X1 U884 ( .IN1(n7014), .IN2(n6634), .IN3(\FIFO[109][7] ), .IN4(n6636), 
        .Q(n1050) );
  AO22X1 U885 ( .IN1(n7003), .IN2(n6634), .IN3(\FIFO[109][8] ), .IN4(n6636), 
        .Q(n1051) );
  AO22X1 U886 ( .IN1(n6992), .IN2(n6634), .IN3(\FIFO[109][9] ), .IN4(n6636), 
        .Q(n1052) );
  AO22X1 U887 ( .IN1(n6981), .IN2(n6634), .IN3(\FIFO[109][10] ), .IN4(n6636), 
        .Q(n1053) );
  AO22X1 U888 ( .IN1(n6970), .IN2(n6634), .IN3(\FIFO[109][11] ), .IN4(n6636), 
        .Q(n1054) );
  AO22X1 U889 ( .IN1(n6959), .IN2(n6634), .IN3(\FIFO[109][12] ), .IN4(n6637), 
        .Q(n1055) );
  AO22X1 U890 ( .IN1(n6948), .IN2(n6634), .IN3(\FIFO[109][13] ), .IN4(n6637), 
        .Q(n1056) );
  AO22X1 U891 ( .IN1(n6937), .IN2(n6633), .IN3(\FIFO[109][14] ), .IN4(n6637), 
        .Q(n1057) );
  AO22X1 U892 ( .IN1(n6926), .IN2(n6633), .IN3(\FIFO[109][15] ), .IN4(n6637), 
        .Q(n1058) );
  AO22X1 U893 ( .IN1(n6915), .IN2(n6633), .IN3(\FIFO[109][16] ), .IN4(n6637), 
        .Q(n1059) );
  AO22X1 U894 ( .IN1(n6904), .IN2(n6633), .IN3(\FIFO[109][17] ), .IN4(n6637), 
        .Q(n1060) );
  AO22X1 U895 ( .IN1(n6893), .IN2(n6633), .IN3(\FIFO[109][18] ), .IN4(n6637), 
        .Q(n1061) );
  AO22X1 U896 ( .IN1(n6882), .IN2(n6633), .IN3(\FIFO[109][19] ), .IN4(n6637), 
        .Q(n1062) );
  AO22X1 U897 ( .IN1(n6871), .IN2(n6633), .IN3(\FIFO[109][20] ), .IN4(n6637), 
        .Q(n1063) );
  AO22X1 U898 ( .IN1(n6860), .IN2(n6635), .IN3(\FIFO[109][21] ), .IN4(n6637), 
        .Q(n1064) );
  AO22X1 U899 ( .IN1(n6849), .IN2(n6634), .IN3(\FIFO[109][22] ), .IN4(n6637), 
        .Q(n1065) );
  AO22X1 U900 ( .IN1(n6838), .IN2(n6633), .IN3(\FIFO[109][23] ), .IN4(n6637), 
        .Q(n1066) );
  AO22X1 U901 ( .IN1(n6827), .IN2(n274), .IN3(\FIFO[109][24] ), .IN4(n6638), 
        .Q(n1067) );
  AO22X1 U902 ( .IN1(n6816), .IN2(n274), .IN3(\FIFO[109][25] ), .IN4(n6638), 
        .Q(n1068) );
  AO22X1 U903 ( .IN1(n6805), .IN2(n274), .IN3(\FIFO[109][26] ), .IN4(n6638), 
        .Q(n1069) );
  AO22X1 U904 ( .IN1(n6794), .IN2(n6635), .IN3(\FIFO[109][27] ), .IN4(n6638), 
        .Q(n1070) );
  AO22X1 U905 ( .IN1(n6783), .IN2(n6635), .IN3(\FIFO[109][28] ), .IN4(n6638), 
        .Q(n1071) );
  AO22X1 U906 ( .IN1(n6772), .IN2(n6634), .IN3(\FIFO[109][29] ), .IN4(n6638), 
        .Q(n1072) );
  AO22X1 U907 ( .IN1(n6761), .IN2(n6633), .IN3(\FIFO[109][30] ), .IN4(n6638), 
        .Q(n1073) );
  AO22X1 U908 ( .IN1(n6750), .IN2(n6634), .IN3(\FIFO[109][31] ), .IN4(n6638), 
        .Q(n1074) );
  AO21X1 U909 ( .IN1(n272), .IN2(n243), .IN3(n5974), .Q(n274) );
  AO22X1 U910 ( .IN1(n7097), .IN2(n6629), .IN3(\FIFO[108][0] ), .IN4(n6630), 
        .Q(n1075) );
  AO22X1 U911 ( .IN1(n7080), .IN2(n6629), .IN3(\FIFO[108][1] ), .IN4(n6630), 
        .Q(n1076) );
  AO22X1 U912 ( .IN1(n7069), .IN2(n6629), .IN3(\FIFO[108][2] ), .IN4(n6630), 
        .Q(n1077) );
  AO22X1 U913 ( .IN1(n7058), .IN2(n6629), .IN3(\FIFO[108][3] ), .IN4(n6630), 
        .Q(n1078) );
  AO22X1 U914 ( .IN1(n7047), .IN2(n6629), .IN3(\FIFO[108][4] ), .IN4(n6630), 
        .Q(n1079) );
  AO22X1 U915 ( .IN1(n7036), .IN2(n6629), .IN3(\FIFO[108][5] ), .IN4(n6630), 
        .Q(n1080) );
  AO22X1 U916 ( .IN1(n7025), .IN2(n6629), .IN3(\FIFO[108][6] ), .IN4(n6630), 
        .Q(n1081) );
  AO22X1 U917 ( .IN1(n7014), .IN2(n6628), .IN3(\FIFO[108][7] ), .IN4(n6630), 
        .Q(n1082) );
  AO22X1 U919 ( .IN1(n6992), .IN2(n6628), .IN3(\FIFO[108][9] ), .IN4(n6630), 
        .Q(n1084) );
  AO22X1 U920 ( .IN1(n6981), .IN2(n6628), .IN3(\FIFO[108][10] ), .IN4(n6630), 
        .Q(n1085) );
  AO22X1 U921 ( .IN1(n6970), .IN2(n6628), .IN3(\FIFO[108][11] ), .IN4(n6630), 
        .Q(n1086) );
  AO22X1 U922 ( .IN1(n6959), .IN2(n6628), .IN3(\FIFO[108][12] ), .IN4(n6631), 
        .Q(n1087) );
  AO22X1 U923 ( .IN1(n6948), .IN2(n6628), .IN3(\FIFO[108][13] ), .IN4(n6631), 
        .Q(n1088) );
  AO22X1 U924 ( .IN1(n6937), .IN2(n6629), .IN3(\FIFO[108][14] ), .IN4(n6631), 
        .Q(n1089) );
  AO22X1 U925 ( .IN1(n6926), .IN2(n6628), .IN3(\FIFO[108][15] ), .IN4(n6631), 
        .Q(n1090) );
  AO22X1 U926 ( .IN1(n6915), .IN2(n6627), .IN3(\FIFO[108][16] ), .IN4(n6631), 
        .Q(n1091) );
  AO22X1 U927 ( .IN1(n6904), .IN2(n6629), .IN3(\FIFO[108][17] ), .IN4(n6631), 
        .Q(n1092) );
  AO22X1 U928 ( .IN1(n6893), .IN2(n6628), .IN3(\FIFO[108][18] ), .IN4(n6631), 
        .Q(n1093) );
  AO22X1 U929 ( .IN1(n6882), .IN2(n6627), .IN3(\FIFO[108][19] ), .IN4(n6631), 
        .Q(n1094) );
  AO22X1 U930 ( .IN1(n6871), .IN2(n6629), .IN3(\FIFO[108][20] ), .IN4(n6631), 
        .Q(n1095) );
  AO22X1 U931 ( .IN1(n6860), .IN2(n6627), .IN3(\FIFO[108][21] ), .IN4(n6631), 
        .Q(n1096) );
  AO22X1 U932 ( .IN1(n6849), .IN2(n6627), .IN3(\FIFO[108][22] ), .IN4(n6631), 
        .Q(n1097) );
  AO22X1 U933 ( .IN1(n6838), .IN2(n6627), .IN3(\FIFO[108][23] ), .IN4(n6631), 
        .Q(n1098) );
  AO22X1 U934 ( .IN1(n6827), .IN2(n6627), .IN3(\FIFO[108][24] ), .IN4(n6632), 
        .Q(n1099) );
  AO22X1 U935 ( .IN1(n6816), .IN2(n6627), .IN3(\FIFO[108][25] ), .IN4(n6632), 
        .Q(n1100) );
  AO22X1 U936 ( .IN1(n6805), .IN2(n6627), .IN3(\FIFO[108][26] ), .IN4(n6632), 
        .Q(n1101) );
  AO22X1 U937 ( .IN1(n6794), .IN2(n6627), .IN3(\FIFO[108][27] ), .IN4(n6632), 
        .Q(n1102) );
  AO22X1 U938 ( .IN1(n6783), .IN2(n6627), .IN3(\FIFO[108][28] ), .IN4(n6632), 
        .Q(n1103) );
  AO22X1 U939 ( .IN1(n6772), .IN2(n6628), .IN3(\FIFO[108][29] ), .IN4(n6632), 
        .Q(n1104) );
  AO22X1 U940 ( .IN1(n6761), .IN2(n6627), .IN3(\FIFO[108][30] ), .IN4(n6632), 
        .Q(n1105) );
  AO22X1 U941 ( .IN1(n6750), .IN2(n6628), .IN3(\FIFO[108][31] ), .IN4(n6632), 
        .Q(n1106) );
  AO21X1 U942 ( .IN1(n272), .IN2(n245), .IN3(n5975), .Q(n275) );
  AO22X1 U967 ( .IN1(n6826), .IN2(n6621), .IN3(\FIFO[107][24] ), .IN4(n6626), 
        .Q(n1131) );
  AO22X1 U968 ( .IN1(n6815), .IN2(n6621), .IN3(\FIFO[107][25] ), .IN4(n6626), 
        .Q(n1132) );
  AO22X1 U969 ( .IN1(n6804), .IN2(n6621), .IN3(\FIFO[107][26] ), .IN4(n6626), 
        .Q(n1133) );
  AO22X1 U970 ( .IN1(n6793), .IN2(n6621), .IN3(\FIFO[107][27] ), .IN4(n6626), 
        .Q(n1134) );
  AO22X1 U971 ( .IN1(n6782), .IN2(n6621), .IN3(\FIFO[107][28] ), .IN4(n6626), 
        .Q(n1135) );
  AO22X1 U972 ( .IN1(n6771), .IN2(n6622), .IN3(\FIFO[107][29] ), .IN4(n6626), 
        .Q(n1136) );
  AO22X1 U973 ( .IN1(n6760), .IN2(n6621), .IN3(\FIFO[107][30] ), .IN4(n6626), 
        .Q(n1137) );
  AO22X1 U974 ( .IN1(n6749), .IN2(n6622), .IN3(\FIFO[107][31] ), .IN4(n6626), 
        .Q(n1138) );
  AO21X1 U975 ( .IN1(n272), .IN2(n247), .IN3(n5974), .Q(n276) );
  AO22X1 U1000 ( .IN1(n6826), .IN2(n277), .IN3(\FIFO[106][24] ), .IN4(n6620), 
        .Q(n1163) );
  AO22X1 U1001 ( .IN1(n6815), .IN2(n277), .IN3(\FIFO[106][25] ), .IN4(n6620), 
        .Q(n1164) );
  AO22X1 U1002 ( .IN1(n6804), .IN2(n277), .IN3(\FIFO[106][26] ), .IN4(n6620), 
        .Q(n1165) );
  AO22X1 U1003 ( .IN1(n6793), .IN2(n6617), .IN3(\FIFO[106][27] ), .IN4(n6620), 
        .Q(n1166) );
  AO22X1 U1004 ( .IN1(n6782), .IN2(n6616), .IN3(\FIFO[106][28] ), .IN4(n6620), 
        .Q(n1167) );
  AO22X1 U1005 ( .IN1(n6771), .IN2(n6617), .IN3(\FIFO[106][29] ), .IN4(n6620), 
        .Q(n1168) );
  AO22X1 U1006 ( .IN1(n6760), .IN2(n6616), .IN3(\FIFO[106][30] ), .IN4(n6620), 
        .Q(n1169) );
  AO22X1 U1007 ( .IN1(n6749), .IN2(n6615), .IN3(\FIFO[106][31] ), .IN4(n6620), 
        .Q(n1170) );
  AO21X1 U1008 ( .IN1(n272), .IN2(n249), .IN3(n5975), .Q(n277) );
  AO22X1 U1009 ( .IN1(n7096), .IN2(n6611), .IN3(\FIFO[105][0] ), .IN4(n6612), 
        .Q(n1171) );
  AO22X1 U1010 ( .IN1(n7079), .IN2(n6611), .IN3(\FIFO[105][1] ), .IN4(n6612), 
        .Q(n1172) );
  AO22X1 U1011 ( .IN1(n7068), .IN2(n6611), .IN3(\FIFO[105][2] ), .IN4(n6612), 
        .Q(n1173) );
  AO22X1 U1012 ( .IN1(n7057), .IN2(n6611), .IN3(\FIFO[105][3] ), .IN4(n6612), 
        .Q(n1174) );
  AO22X1 U1013 ( .IN1(n7046), .IN2(n6611), .IN3(\FIFO[105][4] ), .IN4(n6612), 
        .Q(n1175) );
  AO22X1 U1014 ( .IN1(n7035), .IN2(n6611), .IN3(\FIFO[105][5] ), .IN4(n6612), 
        .Q(n1176) );
  AO22X1 U1015 ( .IN1(n7024), .IN2(n6611), .IN3(\FIFO[105][6] ), .IN4(n6612), 
        .Q(n1177) );
  AO22X1 U1016 ( .IN1(n7013), .IN2(n6610), .IN3(\FIFO[105][7] ), .IN4(n6612), 
        .Q(n1178) );
  AO22X1 U1017 ( .IN1(n7002), .IN2(n6610), .IN3(\FIFO[105][8] ), .IN4(n6612), 
        .Q(n1179) );
  AO22X1 U1018 ( .IN1(n6991), .IN2(n6610), .IN3(\FIFO[105][9] ), .IN4(n6612), 
        .Q(n1180) );
  AO22X1 U1019 ( .IN1(n6980), .IN2(n6610), .IN3(\FIFO[105][10] ), .IN4(n6612), 
        .Q(n1181) );
  AO22X1 U1020 ( .IN1(n6969), .IN2(n6610), .IN3(\FIFO[105][11] ), .IN4(n6612), 
        .Q(n1182) );
  AO22X1 U1021 ( .IN1(n6958), .IN2(n6610), .IN3(\FIFO[105][12] ), .IN4(n6613), 
        .Q(n1183) );
  AO22X1 U1022 ( .IN1(n6947), .IN2(n6610), .IN3(\FIFO[105][13] ), .IN4(n6613), 
        .Q(n1184) );
  AO22X1 U1023 ( .IN1(n6936), .IN2(n6609), .IN3(\FIFO[105][14] ), .IN4(n6613), 
        .Q(n1185) );
  AO22X1 U1024 ( .IN1(n6925), .IN2(n6609), .IN3(\FIFO[105][15] ), .IN4(n6613), 
        .Q(n1186) );
  AO22X1 U1025 ( .IN1(n6914), .IN2(n6609), .IN3(\FIFO[105][16] ), .IN4(n6613), 
        .Q(n1187) );
  AO22X1 U1026 ( .IN1(n6903), .IN2(n6609), .IN3(\FIFO[105][17] ), .IN4(n6613), 
        .Q(n1188) );
  AO22X1 U1027 ( .IN1(n6892), .IN2(n6609), .IN3(\FIFO[105][18] ), .IN4(n6613), 
        .Q(n1189) );
  AO22X1 U1028 ( .IN1(n6881), .IN2(n6609), .IN3(\FIFO[105][19] ), .IN4(n6613), 
        .Q(n1190) );
  AO22X1 U1029 ( .IN1(n6870), .IN2(n6609), .IN3(\FIFO[105][20] ), .IN4(n6613), 
        .Q(n1191) );
  AO22X1 U1030 ( .IN1(n6859), .IN2(n6611), .IN3(\FIFO[105][21] ), .IN4(n6613), 
        .Q(n1192) );
  AO22X1 U1031 ( .IN1(n6848), .IN2(n6610), .IN3(\FIFO[105][22] ), .IN4(n6613), 
        .Q(n1193) );
  AO22X1 U1032 ( .IN1(n6837), .IN2(n6609), .IN3(\FIFO[105][23] ), .IN4(n6613), 
        .Q(n1194) );
  AO22X1 U1033 ( .IN1(n6826), .IN2(n278), .IN3(\FIFO[105][24] ), .IN4(n6614), 
        .Q(n1195) );
  AO22X1 U1034 ( .IN1(n6815), .IN2(n278), .IN3(\FIFO[105][25] ), .IN4(n6614), 
        .Q(n1196) );
  AO22X1 U1035 ( .IN1(n6804), .IN2(n278), .IN3(\FIFO[105][26] ), .IN4(n6614), 
        .Q(n1197) );
  AO22X1 U1036 ( .IN1(n6793), .IN2(n6611), .IN3(\FIFO[105][27] ), .IN4(n6614), 
        .Q(n1198) );
  AO22X1 U1037 ( .IN1(n6782), .IN2(n6610), .IN3(\FIFO[105][28] ), .IN4(n6614), 
        .Q(n1199) );
  AO22X1 U1038 ( .IN1(n6771), .IN2(n6611), .IN3(\FIFO[105][29] ), .IN4(n6614), 
        .Q(n1200) );
  AO22X1 U1039 ( .IN1(n6760), .IN2(n6610), .IN3(\FIFO[105][30] ), .IN4(n6614), 
        .Q(n1201) );
  AO22X1 U1040 ( .IN1(n6749), .IN2(n6609), .IN3(\FIFO[105][31] ), .IN4(n6614), 
        .Q(n1202) );
  AO21X1 U1041 ( .IN1(n272), .IN2(n251), .IN3(n5974), .Q(n278) );
  AO22X1 U1042 ( .IN1(n7096), .IN2(n6605), .IN3(\FIFO[104][0] ), .IN4(n6606), 
        .Q(n1203) );
  AO22X1 U1043 ( .IN1(n7079), .IN2(n6605), .IN3(\FIFO[104][1] ), .IN4(n6606), 
        .Q(n1204) );
  AO22X1 U1044 ( .IN1(n7068), .IN2(n6605), .IN3(\FIFO[104][2] ), .IN4(n6606), 
        .Q(n1205) );
  AO22X1 U1045 ( .IN1(n7057), .IN2(n6605), .IN3(\FIFO[104][3] ), .IN4(n6606), 
        .Q(n1206) );
  AO22X1 U1046 ( .IN1(n7046), .IN2(n6605), .IN3(\FIFO[104][4] ), .IN4(n6606), 
        .Q(n1207) );
  AO22X1 U1047 ( .IN1(n7035), .IN2(n6605), .IN3(\FIFO[104][5] ), .IN4(n6606), 
        .Q(n1208) );
  AO22X1 U1048 ( .IN1(n7024), .IN2(n6605), .IN3(\FIFO[104][6] ), .IN4(n6606), 
        .Q(n1209) );
  AO22X1 U1049 ( .IN1(n7013), .IN2(n6604), .IN3(\FIFO[104][7] ), .IN4(n6606), 
        .Q(n1210) );
  AO22X1 U1050 ( .IN1(n7002), .IN2(n6604), .IN3(\FIFO[104][8] ), .IN4(n6606), 
        .Q(n1211) );
  AO22X1 U1051 ( .IN1(n6991), .IN2(n6604), .IN3(\FIFO[104][9] ), .IN4(n6606), 
        .Q(n1212) );
  AO22X1 U1052 ( .IN1(n6980), .IN2(n6604), .IN3(\FIFO[104][10] ), .IN4(n6606), 
        .Q(n1213) );
  AO22X1 U1053 ( .IN1(n6969), .IN2(n6604), .IN3(\FIFO[104][11] ), .IN4(n6606), 
        .Q(n1214) );
  AO22X1 U1054 ( .IN1(n6958), .IN2(n6604), .IN3(\FIFO[104][12] ), .IN4(n6607), 
        .Q(n1215) );
  AO22X1 U1055 ( .IN1(n6947), .IN2(n6604), .IN3(\FIFO[104][13] ), .IN4(n6607), 
        .Q(n1216) );
  AO22X1 U1056 ( .IN1(n6936), .IN2(n6603), .IN3(\FIFO[104][14] ), .IN4(n6607), 
        .Q(n1217) );
  AO22X1 U1057 ( .IN1(n6925), .IN2(n6603), .IN3(\FIFO[104][15] ), .IN4(n6607), 
        .Q(n1218) );
  AO22X1 U1058 ( .IN1(n6914), .IN2(n6603), .IN3(\FIFO[104][16] ), .IN4(n6607), 
        .Q(n1219) );
  AO22X1 U1059 ( .IN1(n6903), .IN2(n6603), .IN3(\FIFO[104][17] ), .IN4(n6607), 
        .Q(n1220) );
  AO22X1 U1060 ( .IN1(n6892), .IN2(n6603), .IN3(\FIFO[104][18] ), .IN4(n6607), 
        .Q(n1221) );
  AO22X1 U1061 ( .IN1(n6881), .IN2(n6603), .IN3(\FIFO[104][19] ), .IN4(n6607), 
        .Q(n1222) );
  AO22X1 U1062 ( .IN1(n6870), .IN2(n6603), .IN3(\FIFO[104][20] ), .IN4(n6607), 
        .Q(n1223) );
  AO22X1 U1063 ( .IN1(n6859), .IN2(n6605), .IN3(\FIFO[104][21] ), .IN4(n6607), 
        .Q(n1224) );
  AO22X1 U1064 ( .IN1(n6848), .IN2(n6604), .IN3(\FIFO[104][22] ), .IN4(n6607), 
        .Q(n1225) );
  AO22X1 U1065 ( .IN1(n6837), .IN2(n6603), .IN3(\FIFO[104][23] ), .IN4(n6607), 
        .Q(n1226) );
  AO22X1 U1066 ( .IN1(n6826), .IN2(n279), .IN3(\FIFO[104][24] ), .IN4(n6608), 
        .Q(n1227) );
  AO22X1 U1067 ( .IN1(n6815), .IN2(n279), .IN3(\FIFO[104][25] ), .IN4(n6608), 
        .Q(n1228) );
  AO22X1 U1068 ( .IN1(n6804), .IN2(n279), .IN3(\FIFO[104][26] ), .IN4(n6608), 
        .Q(n1229) );
  AO22X1 U1069 ( .IN1(n6793), .IN2(n6605), .IN3(\FIFO[104][27] ), .IN4(n6608), 
        .Q(n1230) );
  AO22X1 U1070 ( .IN1(n6782), .IN2(n6605), .IN3(\FIFO[104][28] ), .IN4(n6608), 
        .Q(n1231) );
  AO22X1 U1071 ( .IN1(n6771), .IN2(n6604), .IN3(\FIFO[104][29] ), .IN4(n6608), 
        .Q(n1232) );
  AO22X1 U1072 ( .IN1(n6760), .IN2(n6603), .IN3(\FIFO[104][30] ), .IN4(n6608), 
        .Q(n1233) );
  AO22X1 U1073 ( .IN1(n6749), .IN2(n6604), .IN3(\FIFO[104][31] ), .IN4(n6608), 
        .Q(n1234) );
  AO21X1 U1074 ( .IN1(n272), .IN2(n253), .IN3(n5975), .Q(n279) );
  AO22X1 U1099 ( .IN1(n6826), .IN2(n6597), .IN3(\FIFO[103][24] ), .IN4(n6602), 
        .Q(n1259) );
  AO22X1 U1100 ( .IN1(n6815), .IN2(n6597), .IN3(\FIFO[103][25] ), .IN4(n6602), 
        .Q(n1260) );
  AO22X1 U1101 ( .IN1(n6804), .IN2(n6597), .IN3(\FIFO[103][26] ), .IN4(n6602), 
        .Q(n1261) );
  AO22X1 U1102 ( .IN1(n6793), .IN2(n6597), .IN3(\FIFO[103][27] ), .IN4(n6602), 
        .Q(n1262) );
  AO22X1 U1103 ( .IN1(n6782), .IN2(n6597), .IN3(\FIFO[103][28] ), .IN4(n6602), 
        .Q(n1263) );
  AO22X1 U1104 ( .IN1(n6771), .IN2(n6598), .IN3(\FIFO[103][29] ), .IN4(n6602), 
        .Q(n1264) );
  AO22X1 U1105 ( .IN1(n6760), .IN2(n6597), .IN3(\FIFO[103][30] ), .IN4(n6602), 
        .Q(n1265) );
  AO22X1 U1106 ( .IN1(n6749), .IN2(n6598), .IN3(\FIFO[103][31] ), .IN4(n6602), 
        .Q(n1266) );
  AO21X1 U1107 ( .IN1(n272), .IN2(n255), .IN3(n5974), .Q(n280) );
  AO22X1 U1132 ( .IN1(n6826), .IN2(n6591), .IN3(\FIFO[102][24] ), .IN4(n6596), 
        .Q(n1291) );
  AO22X1 U1133 ( .IN1(n6815), .IN2(n6591), .IN3(\FIFO[102][25] ), .IN4(n6596), 
        .Q(n1292) );
  AO22X1 U1134 ( .IN1(n6804), .IN2(n6591), .IN3(\FIFO[102][26] ), .IN4(n6596), 
        .Q(n1293) );
  AO22X1 U1135 ( .IN1(n6793), .IN2(n6591), .IN3(\FIFO[102][27] ), .IN4(n6596), 
        .Q(n1294) );
  AO22X1 U1136 ( .IN1(n6782), .IN2(n6591), .IN3(\FIFO[102][28] ), .IN4(n6596), 
        .Q(n1295) );
  AO22X1 U1137 ( .IN1(n6771), .IN2(n6592), .IN3(\FIFO[102][29] ), .IN4(n6596), 
        .Q(n1296) );
  AO22X1 U1138 ( .IN1(n6760), .IN2(n6591), .IN3(\FIFO[102][30] ), .IN4(n6596), 
        .Q(n1297) );
  AO22X1 U1139 ( .IN1(n6749), .IN2(n6592), .IN3(\FIFO[102][31] ), .IN4(n6596), 
        .Q(n1298) );
  AO21X1 U1140 ( .IN1(n272), .IN2(n257), .IN3(n5975), .Q(n281) );
  AO22X1 U1141 ( .IN1(n7096), .IN2(n6587), .IN3(\FIFO[101][0] ), .IN4(n6588), 
        .Q(n1299) );
  AO22X1 U1142 ( .IN1(n7079), .IN2(n6587), .IN3(\FIFO[101][1] ), .IN4(n6588), 
        .Q(n1300) );
  AO22X1 U1143 ( .IN1(n7068), .IN2(n6587), .IN3(\FIFO[101][2] ), .IN4(n6588), 
        .Q(n1301) );
  AO22X1 U1144 ( .IN1(n7057), .IN2(n6587), .IN3(\FIFO[101][3] ), .IN4(n6588), 
        .Q(n1302) );
  AO22X1 U1145 ( .IN1(n7046), .IN2(n6587), .IN3(\FIFO[101][4] ), .IN4(n6588), 
        .Q(n1303) );
  AO22X1 U1146 ( .IN1(n7035), .IN2(n6587), .IN3(\FIFO[101][5] ), .IN4(n6588), 
        .Q(n1304) );
  AO22X1 U1147 ( .IN1(n7024), .IN2(n6587), .IN3(\FIFO[101][6] ), .IN4(n6588), 
        .Q(n1305) );
  AO22X1 U1148 ( .IN1(n7013), .IN2(n6586), .IN3(\FIFO[101][7] ), .IN4(n6588), 
        .Q(n1306) );
  AO22X1 U1149 ( .IN1(n7002), .IN2(n6586), .IN3(\FIFO[101][8] ), .IN4(n6588), 
        .Q(n1307) );
  AO22X1 U1150 ( .IN1(n6991), .IN2(n6586), .IN3(\FIFO[101][9] ), .IN4(n6588), 
        .Q(n1308) );
  AO22X1 U1151 ( .IN1(n6980), .IN2(n6586), .IN3(\FIFO[101][10] ), .IN4(n6588), 
        .Q(n1309) );
  AO22X1 U1152 ( .IN1(n6969), .IN2(n6586), .IN3(\FIFO[101][11] ), .IN4(n6588), 
        .Q(n1310) );
  AO22X1 U1153 ( .IN1(n6958), .IN2(n6586), .IN3(\FIFO[101][12] ), .IN4(n6589), 
        .Q(n1311) );
  AO22X1 U1154 ( .IN1(n6947), .IN2(n6586), .IN3(\FIFO[101][13] ), .IN4(n6589), 
        .Q(n1312) );
  AO22X1 U1155 ( .IN1(n6936), .IN2(n6585), .IN3(\FIFO[101][14] ), .IN4(n6589), 
        .Q(n1313) );
  AO22X1 U1156 ( .IN1(n6925), .IN2(n6585), .IN3(\FIFO[101][15] ), .IN4(n6589), 
        .Q(n1314) );
  AO22X1 U1157 ( .IN1(n6914), .IN2(n6585), .IN3(\FIFO[101][16] ), .IN4(n6589), 
        .Q(n1315) );
  AO22X1 U1158 ( .IN1(n6903), .IN2(n6585), .IN3(\FIFO[101][17] ), .IN4(n6589), 
        .Q(n1316) );
  AO22X1 U1159 ( .IN1(n6892), .IN2(n6585), .IN3(\FIFO[101][18] ), .IN4(n6589), 
        .Q(n1317) );
  AO22X1 U1160 ( .IN1(n6881), .IN2(n6585), .IN3(\FIFO[101][19] ), .IN4(n6589), 
        .Q(n1318) );
  AO22X1 U1161 ( .IN1(n6870), .IN2(n6585), .IN3(\FIFO[101][20] ), .IN4(n6589), 
        .Q(n1319) );
  AO22X1 U1162 ( .IN1(n6859), .IN2(n6587), .IN3(\FIFO[101][21] ), .IN4(n6589), 
        .Q(n1320) );
  AO22X1 U1163 ( .IN1(n6848), .IN2(n6586), .IN3(\FIFO[101][22] ), .IN4(n6589), 
        .Q(n1321) );
  AO22X1 U1164 ( .IN1(n6837), .IN2(n6585), .IN3(\FIFO[101][23] ), .IN4(n6589), 
        .Q(n1322) );
  AO22X1 U1165 ( .IN1(n6826), .IN2(n282), .IN3(\FIFO[101][24] ), .IN4(n6590), 
        .Q(n1323) );
  AO22X1 U1166 ( .IN1(n6815), .IN2(n282), .IN3(\FIFO[101][25] ), .IN4(n6590), 
        .Q(n1324) );
  AO22X1 U1167 ( .IN1(n6804), .IN2(n282), .IN3(\FIFO[101][26] ), .IN4(n6590), 
        .Q(n1325) );
  AO22X1 U1168 ( .IN1(n6793), .IN2(n6587), .IN3(\FIFO[101][27] ), .IN4(n6590), 
        .Q(n1326) );
  AO22X1 U1169 ( .IN1(n6782), .IN2(n6586), .IN3(\FIFO[101][28] ), .IN4(n6590), 
        .Q(n1327) );
  AO22X1 U1170 ( .IN1(n6771), .IN2(n6587), .IN3(\FIFO[101][29] ), .IN4(n6590), 
        .Q(n1328) );
  AO22X1 U1171 ( .IN1(n6760), .IN2(n6586), .IN3(\FIFO[101][30] ), .IN4(n6590), 
        .Q(n1329) );
  AO22X1 U1172 ( .IN1(n6749), .IN2(n6585), .IN3(\FIFO[101][31] ), .IN4(n6590), 
        .Q(n1330) );
  AO21X1 U1173 ( .IN1(n272), .IN2(n259), .IN3(n5974), .Q(n282) );
  AO22X1 U1174 ( .IN1(n7096), .IN2(n6581), .IN3(\FIFO[100][0] ), .IN4(n6582), 
        .Q(n1331) );
  AO22X1 U1175 ( .IN1(n7079), .IN2(n6581), .IN3(\FIFO[100][1] ), .IN4(n6582), 
        .Q(n1332) );
  AO22X1 U1176 ( .IN1(n7068), .IN2(n6581), .IN3(\FIFO[100][2] ), .IN4(n6582), 
        .Q(n1333) );
  AO22X1 U1177 ( .IN1(n7057), .IN2(n6581), .IN3(\FIFO[100][3] ), .IN4(n6582), 
        .Q(n1334) );
  AO22X1 U1178 ( .IN1(n7046), .IN2(n6581), .IN3(\FIFO[100][4] ), .IN4(n6582), 
        .Q(n1335) );
  AO22X1 U1179 ( .IN1(n7035), .IN2(n6581), .IN3(\FIFO[100][5] ), .IN4(n6582), 
        .Q(n1336) );
  AO22X1 U1180 ( .IN1(n7024), .IN2(n6581), .IN3(\FIFO[100][6] ), .IN4(n6582), 
        .Q(n1337) );
  AO22X1 U1181 ( .IN1(n7013), .IN2(n6580), .IN3(\FIFO[100][7] ), .IN4(n6582), 
        .Q(n1338) );
  AO22X1 U1182 ( .IN1(n7002), .IN2(n6580), .IN3(\FIFO[100][8] ), .IN4(n6582), 
        .Q(n1339) );
  AO22X1 U1183 ( .IN1(n6991), .IN2(n6580), .IN3(\FIFO[100][9] ), .IN4(n6582), 
        .Q(n1340) );
  AO22X1 U1184 ( .IN1(n6980), .IN2(n6580), .IN3(\FIFO[100][10] ), .IN4(n6582), 
        .Q(n1341) );
  AO22X1 U1185 ( .IN1(n6969), .IN2(n6580), .IN3(\FIFO[100][11] ), .IN4(n6582), 
        .Q(n1342) );
  AO22X1 U1186 ( .IN1(n6958), .IN2(n6580), .IN3(\FIFO[100][12] ), .IN4(n6583), 
        .Q(n1343) );
  AO22X1 U1187 ( .IN1(n6947), .IN2(n6580), .IN3(\FIFO[100][13] ), .IN4(n6583), 
        .Q(n1344) );
  AO22X1 U1188 ( .IN1(n6936), .IN2(n6579), .IN3(\FIFO[100][14] ), .IN4(n6583), 
        .Q(n1345) );
  AO22X1 U1189 ( .IN1(n6925), .IN2(n6579), .IN3(\FIFO[100][15] ), .IN4(n6583), 
        .Q(n1346) );
  AO22X1 U1190 ( .IN1(n6914), .IN2(n6579), .IN3(\FIFO[100][16] ), .IN4(n6583), 
        .Q(n1347) );
  AO22X1 U1191 ( .IN1(n6903), .IN2(n6579), .IN3(\FIFO[100][17] ), .IN4(n6583), 
        .Q(n1348) );
  AO22X1 U1192 ( .IN1(n6892), .IN2(n6579), .IN3(\FIFO[100][18] ), .IN4(n6583), 
        .Q(n1349) );
  AO22X1 U1193 ( .IN1(n6881), .IN2(n6579), .IN3(\FIFO[100][19] ), .IN4(n6583), 
        .Q(n1350) );
  AO22X1 U1194 ( .IN1(n6870), .IN2(n6579), .IN3(\FIFO[100][20] ), .IN4(n6583), 
        .Q(n1351) );
  AO22X1 U1195 ( .IN1(n6859), .IN2(n6581), .IN3(\FIFO[100][21] ), .IN4(n6583), 
        .Q(n1352) );
  AO22X1 U1196 ( .IN1(n6848), .IN2(n6580), .IN3(\FIFO[100][22] ), .IN4(n6583), 
        .Q(n1353) );
  AO22X1 U1197 ( .IN1(n6837), .IN2(n6579), .IN3(\FIFO[100][23] ), .IN4(n6583), 
        .Q(n1354) );
  AO22X1 U1198 ( .IN1(n6826), .IN2(n283), .IN3(\FIFO[100][24] ), .IN4(n6584), 
        .Q(n1355) );
  AO22X1 U1199 ( .IN1(n6815), .IN2(n283), .IN3(\FIFO[100][25] ), .IN4(n6584), 
        .Q(n1356) );
  AO22X1 U1200 ( .IN1(n6804), .IN2(n283), .IN3(\FIFO[100][26] ), .IN4(n6584), 
        .Q(n1357) );
  AO22X1 U1201 ( .IN1(n6793), .IN2(n6581), .IN3(\FIFO[100][27] ), .IN4(n6584), 
        .Q(n1358) );
  AO22X1 U1202 ( .IN1(n6782), .IN2(n6580), .IN3(\FIFO[100][28] ), .IN4(n6584), 
        .Q(n1359) );
  AO22X1 U1203 ( .IN1(n6771), .IN2(n6581), .IN3(\FIFO[100][29] ), .IN4(n6584), 
        .Q(n1360) );
  AO22X1 U1204 ( .IN1(n6760), .IN2(n6580), .IN3(\FIFO[100][30] ), .IN4(n6584), 
        .Q(n1361) );
  AO22X1 U1205 ( .IN1(n6749), .IN2(n6579), .IN3(\FIFO[100][31] ), .IN4(n6584), 
        .Q(n1362) );
  AO21X1 U1206 ( .IN1(n272), .IN2(n261), .IN3(n5975), .Q(n283) );
  AO22X1 U1231 ( .IN1(n6826), .IN2(n284), .IN3(\FIFO[99][24] ), .IN4(n6578), 
        .Q(n1387) );
  AO22X1 U1232 ( .IN1(n6815), .IN2(n284), .IN3(\FIFO[99][25] ), .IN4(n6578), 
        .Q(n1388) );
  AO22X1 U1233 ( .IN1(n6804), .IN2(n284), .IN3(\FIFO[99][26] ), .IN4(n6578), 
        .Q(n1389) );
  AO22X1 U1234 ( .IN1(n6793), .IN2(n6575), .IN3(\FIFO[99][27] ), .IN4(n6578), 
        .Q(n1390) );
  AO22X1 U1235 ( .IN1(n6782), .IN2(n6575), .IN3(\FIFO[99][28] ), .IN4(n6578), 
        .Q(n1391) );
  AO22X1 U1236 ( .IN1(n6771), .IN2(n6574), .IN3(\FIFO[99][29] ), .IN4(n6578), 
        .Q(n1392) );
  AO22X1 U1237 ( .IN1(n6760), .IN2(n6573), .IN3(\FIFO[99][30] ), .IN4(n6578), 
        .Q(n1393) );
  AO22X1 U1238 ( .IN1(n6749), .IN2(n6574), .IN3(\FIFO[99][31] ), .IN4(n6578), 
        .Q(n1394) );
  AO21X1 U1239 ( .IN1(n272), .IN2(n263), .IN3(n5974), .Q(n284) );
  AO22X1 U1264 ( .IN1(n6826), .IN2(n6567), .IN3(\FIFO[98][24] ), .IN4(n6572), 
        .Q(n1419) );
  AO22X1 U1265 ( .IN1(n6815), .IN2(n6567), .IN3(\FIFO[98][25] ), .IN4(n6572), 
        .Q(n1420) );
  AO22X1 U1266 ( .IN1(n6804), .IN2(n6567), .IN3(\FIFO[98][26] ), .IN4(n6572), 
        .Q(n1421) );
  AO22X1 U1267 ( .IN1(n6793), .IN2(n6567), .IN3(\FIFO[98][27] ), .IN4(n6572), 
        .Q(n1422) );
  AO22X1 U1268 ( .IN1(n6782), .IN2(n6567), .IN3(\FIFO[98][28] ), .IN4(n6572), 
        .Q(n1423) );
  AO22X1 U1269 ( .IN1(n6771), .IN2(n6568), .IN3(\FIFO[98][29] ), .IN4(n6572), 
        .Q(n1424) );
  AO22X1 U1270 ( .IN1(n6760), .IN2(n6567), .IN3(\FIFO[98][30] ), .IN4(n6572), 
        .Q(n1425) );
  AO22X1 U1271 ( .IN1(n6749), .IN2(n6568), .IN3(\FIFO[98][31] ), .IN4(n6572), 
        .Q(n1426) );
  AO21X1 U1272 ( .IN1(n272), .IN2(n265), .IN3(n5975), .Q(n285) );
  AO22X1 U1274 ( .IN1(n7079), .IN2(n6562), .IN3(\FIFO[97][1] ), .IN4(n6564), 
        .Q(n1428) );
  AO22X1 U1275 ( .IN1(n7068), .IN2(n6561), .IN3(\FIFO[97][2] ), .IN4(n6564), 
        .Q(n1429) );
  AO22X1 U1276 ( .IN1(n7057), .IN2(n6563), .IN3(\FIFO[97][3] ), .IN4(n6564), 
        .Q(n1430) );
  AO22X1 U1277 ( .IN1(n7046), .IN2(n6562), .IN3(\FIFO[97][4] ), .IN4(n6564), 
        .Q(n1431) );
  AO22X1 U1278 ( .IN1(n7035), .IN2(n6561), .IN3(\FIFO[97][5] ), .IN4(n6564), 
        .Q(n1432) );
  AO22X1 U1279 ( .IN1(n7024), .IN2(n6563), .IN3(\FIFO[97][6] ), .IN4(n6564), 
        .Q(n1433) );
  AO22X1 U1280 ( .IN1(n7013), .IN2(n6563), .IN3(\FIFO[97][7] ), .IN4(n6564), 
        .Q(n1434) );
  AO22X1 U1281 ( .IN1(n7002), .IN2(n6563), .IN3(\FIFO[97][8] ), .IN4(n6564), 
        .Q(n1435) );
  AO22X1 U1282 ( .IN1(n6991), .IN2(n6563), .IN3(\FIFO[97][9] ), .IN4(n6564), 
        .Q(n1436) );
  AO22X1 U1283 ( .IN1(n6980), .IN2(n6563), .IN3(\FIFO[97][10] ), .IN4(n6564), 
        .Q(n1437) );
  AO22X1 U1284 ( .IN1(n6969), .IN2(n6563), .IN3(\FIFO[97][11] ), .IN4(n6564), 
        .Q(n1438) );
  AO22X1 U1285 ( .IN1(n6958), .IN2(n6563), .IN3(\FIFO[97][12] ), .IN4(n6565), 
        .Q(n1439) );
  AO22X1 U1286 ( .IN1(n6947), .IN2(n6563), .IN3(\FIFO[97][13] ), .IN4(n6565), 
        .Q(n1440) );
  AO22X1 U1288 ( .IN1(n6925), .IN2(n6562), .IN3(\FIFO[97][15] ), .IN4(n6565), 
        .Q(n1442) );
  AO22X1 U1289 ( .IN1(n6914), .IN2(n6562), .IN3(\FIFO[97][16] ), .IN4(n6565), 
        .Q(n1443) );
  AO22X1 U1290 ( .IN1(n6903), .IN2(n6562), .IN3(\FIFO[97][17] ), .IN4(n6565), 
        .Q(n1444) );
  AO22X1 U1291 ( .IN1(n6892), .IN2(n6562), .IN3(\FIFO[97][18] ), .IN4(n6565), 
        .Q(n1445) );
  AO22X1 U1292 ( .IN1(n6881), .IN2(n6562), .IN3(\FIFO[97][19] ), .IN4(n6565), 
        .Q(n1446) );
  AO22X1 U1293 ( .IN1(n6870), .IN2(n6562), .IN3(\FIFO[97][20] ), .IN4(n6565), 
        .Q(n1447) );
  AO22X1 U1294 ( .IN1(n6859), .IN2(n6561), .IN3(\FIFO[97][21] ), .IN4(n6565), 
        .Q(n1448) );
  AO22X1 U1295 ( .IN1(n6848), .IN2(n6561), .IN3(\FIFO[97][22] ), .IN4(n6565), 
        .Q(n1449) );
  AO22X1 U1296 ( .IN1(n6837), .IN2(n6561), .IN3(\FIFO[97][23] ), .IN4(n6565), 
        .Q(n1450) );
  AO22X1 U1297 ( .IN1(n6826), .IN2(n6561), .IN3(\FIFO[97][24] ), .IN4(n6566), 
        .Q(n1451) );
  AO22X1 U1298 ( .IN1(n6815), .IN2(n6561), .IN3(\FIFO[97][25] ), .IN4(n6566), 
        .Q(n1452) );
  AO22X1 U1299 ( .IN1(n6804), .IN2(n6561), .IN3(\FIFO[97][26] ), .IN4(n6566), 
        .Q(n1453) );
  AO22X1 U1300 ( .IN1(n6793), .IN2(n6561), .IN3(\FIFO[97][27] ), .IN4(n6566), 
        .Q(n1454) );
  AO22X1 U1301 ( .IN1(n6782), .IN2(n6561), .IN3(\FIFO[97][28] ), .IN4(n6566), 
        .Q(n1455) );
  AO22X1 U1302 ( .IN1(n6771), .IN2(n6562), .IN3(\FIFO[97][29] ), .IN4(n6566), 
        .Q(n1456) );
  AO22X1 U1303 ( .IN1(n6760), .IN2(n6561), .IN3(\FIFO[97][30] ), .IN4(n6566), 
        .Q(n1457) );
  AO22X1 U1304 ( .IN1(n6749), .IN2(n6562), .IN3(\FIFO[97][31] ), .IN4(n6566), 
        .Q(n1458) );
  AO21X1 U1305 ( .IN1(n272), .IN2(n267), .IN3(n5973), .Q(n286) );
  AO22X1 U1306 ( .IN1(n7096), .IN2(n6557), .IN3(\FIFO[96][0] ), .IN4(n6558), 
        .Q(n1459) );
  AO22X1 U1307 ( .IN1(n7079), .IN2(n6557), .IN3(\FIFO[96][1] ), .IN4(n6558), 
        .Q(n1460) );
  AO22X1 U1308 ( .IN1(n7068), .IN2(n6557), .IN3(\FIFO[96][2] ), .IN4(n6558), 
        .Q(n1461) );
  AO22X1 U1309 ( .IN1(n7057), .IN2(n6557), .IN3(\FIFO[96][3] ), .IN4(n6558), 
        .Q(n1462) );
  AO22X1 U1310 ( .IN1(n7046), .IN2(n6557), .IN3(\FIFO[96][4] ), .IN4(n6558), 
        .Q(n1463) );
  AO22X1 U1311 ( .IN1(n7035), .IN2(n6557), .IN3(\FIFO[96][5] ), .IN4(n6558), 
        .Q(n1464) );
  AO22X1 U1312 ( .IN1(n7024), .IN2(n6557), .IN3(\FIFO[96][6] ), .IN4(n6558), 
        .Q(n1465) );
  AO22X1 U1313 ( .IN1(n7013), .IN2(n6556), .IN3(\FIFO[96][7] ), .IN4(n6558), 
        .Q(n1466) );
  AO22X1 U1314 ( .IN1(n7002), .IN2(n6556), .IN3(\FIFO[96][8] ), .IN4(n6558), 
        .Q(n1467) );
  AO22X1 U1315 ( .IN1(n6991), .IN2(n6556), .IN3(\FIFO[96][9] ), .IN4(n6558), 
        .Q(n1468) );
  AO22X1 U1316 ( .IN1(n6980), .IN2(n6556), .IN3(\FIFO[96][10] ), .IN4(n6558), 
        .Q(n1469) );
  AO22X1 U1317 ( .IN1(n6969), .IN2(n6556), .IN3(\FIFO[96][11] ), .IN4(n6558), 
        .Q(n1470) );
  AO22X1 U1318 ( .IN1(n6958), .IN2(n6556), .IN3(\FIFO[96][12] ), .IN4(n6559), 
        .Q(n1471) );
  AO22X1 U1319 ( .IN1(n6947), .IN2(n6556), .IN3(\FIFO[96][13] ), .IN4(n6559), 
        .Q(n1472) );
  AO22X1 U1320 ( .IN1(n6936), .IN2(n6555), .IN3(\FIFO[96][14] ), .IN4(n6559), 
        .Q(n1473) );
  AO22X1 U1321 ( .IN1(n6925), .IN2(n6555), .IN3(\FIFO[96][15] ), .IN4(n6559), 
        .Q(n1474) );
  AO22X1 U1322 ( .IN1(n6914), .IN2(n6555), .IN3(\FIFO[96][16] ), .IN4(n6559), 
        .Q(n1475) );
  AO22X1 U1323 ( .IN1(n6903), .IN2(n6555), .IN3(\FIFO[96][17] ), .IN4(n6559), 
        .Q(n1476) );
  AO22X1 U1324 ( .IN1(n6892), .IN2(n6555), .IN3(\FIFO[96][18] ), .IN4(n6559), 
        .Q(n1477) );
  AO22X1 U1325 ( .IN1(n6881), .IN2(n6555), .IN3(\FIFO[96][19] ), .IN4(n6559), 
        .Q(n1478) );
  AO22X1 U1326 ( .IN1(n6870), .IN2(n6555), .IN3(\FIFO[96][20] ), .IN4(n6559), 
        .Q(n1479) );
  AO22X1 U1327 ( .IN1(n6859), .IN2(n6557), .IN3(\FIFO[96][21] ), .IN4(n6559), 
        .Q(n1480) );
  AO22X1 U1328 ( .IN1(n6848), .IN2(n6556), .IN3(\FIFO[96][22] ), .IN4(n6559), 
        .Q(n1481) );
  AO22X1 U1329 ( .IN1(n6837), .IN2(n6555), .IN3(\FIFO[96][23] ), .IN4(n6559), 
        .Q(n1482) );
  AO22X1 U1330 ( .IN1(n6826), .IN2(n287), .IN3(\FIFO[96][24] ), .IN4(n6560), 
        .Q(n1483) );
  AO22X1 U1331 ( .IN1(n6815), .IN2(n287), .IN3(\FIFO[96][25] ), .IN4(n6560), 
        .Q(n1484) );
  AO22X1 U1332 ( .IN1(n6804), .IN2(n287), .IN3(\FIFO[96][26] ), .IN4(n6560), 
        .Q(n1485) );
  AO22X1 U1333 ( .IN1(n6793), .IN2(n6557), .IN3(\FIFO[96][27] ), .IN4(n6560), 
        .Q(n1486) );
  AO22X1 U1334 ( .IN1(n6782), .IN2(n6556), .IN3(\FIFO[96][28] ), .IN4(n6560), 
        .Q(n1487) );
  AO22X1 U1335 ( .IN1(n6771), .IN2(n6557), .IN3(\FIFO[96][29] ), .IN4(n6560), 
        .Q(n1488) );
  AO22X1 U1336 ( .IN1(n6760), .IN2(n6556), .IN3(\FIFO[96][30] ), .IN4(n6560), 
        .Q(n1489) );
  AO22X1 U1337 ( .IN1(n6749), .IN2(n6555), .IN3(\FIFO[96][31] ), .IN4(n6560), 
        .Q(n1490) );
  AO21X1 U1338 ( .IN1(n272), .IN2(n269), .IN3(n5973), .Q(n287) );
  AO22X1 U1364 ( .IN1(n6825), .IN2(n288), .IN3(\FIFO[95][24] ), .IN4(n6554), 
        .Q(n1515) );
  AO22X1 U1365 ( .IN1(n6814), .IN2(n288), .IN3(\FIFO[95][25] ), .IN4(n6554), 
        .Q(n1516) );
  AO22X1 U1366 ( .IN1(n6803), .IN2(n288), .IN3(\FIFO[95][26] ), .IN4(n6554), 
        .Q(n1517) );
  AO22X1 U1367 ( .IN1(n6792), .IN2(n6551), .IN3(\FIFO[95][27] ), .IN4(n6554), 
        .Q(n1518) );
  AO22X1 U1368 ( .IN1(n6781), .IN2(n6551), .IN3(\FIFO[95][28] ), .IN4(n6554), 
        .Q(n1519) );
  AO22X1 U1369 ( .IN1(n6770), .IN2(n6550), .IN3(\FIFO[95][29] ), .IN4(n6554), 
        .Q(n1520) );
  AO22X1 U1370 ( .IN1(n6759), .IN2(n6549), .IN3(\FIFO[95][30] ), .IN4(n6554), 
        .Q(n1521) );
  AO22X1 U1371 ( .IN1(n6748), .IN2(n6550), .IN3(\FIFO[95][31] ), .IN4(n6554), 
        .Q(n1522) );
  AO21X1 U1372 ( .IN1(n289), .IN2(n238), .IN3(n5973), .Q(n288) );
  AO22X1 U1397 ( .IN1(n6825), .IN2(n6543), .IN3(\FIFO[94][24] ), .IN4(n6548), 
        .Q(n1547) );
  AO22X1 U1398 ( .IN1(n6814), .IN2(n6543), .IN3(\FIFO[94][25] ), .IN4(n6548), 
        .Q(n1548) );
  AO22X1 U1399 ( .IN1(n6803), .IN2(n6543), .IN3(\FIFO[94][26] ), .IN4(n6548), 
        .Q(n1549) );
  AO22X1 U1400 ( .IN1(n6792), .IN2(n6543), .IN3(\FIFO[94][27] ), .IN4(n6548), 
        .Q(n1550) );
  AO22X1 U1401 ( .IN1(n6781), .IN2(n6543), .IN3(\FIFO[94][28] ), .IN4(n6548), 
        .Q(n1551) );
  AO22X1 U1402 ( .IN1(n6770), .IN2(n6544), .IN3(\FIFO[94][29] ), .IN4(n6548), 
        .Q(n1552) );
  AO22X1 U1403 ( .IN1(n6759), .IN2(n6543), .IN3(\FIFO[94][30] ), .IN4(n6548), 
        .Q(n1553) );
  AO22X1 U1404 ( .IN1(n6748), .IN2(n6544), .IN3(\FIFO[94][31] ), .IN4(n6548), 
        .Q(n1554) );
  AO21X1 U1405 ( .IN1(n289), .IN2(n241), .IN3(n7359), .Q(n290) );
  AO22X1 U1406 ( .IN1(n7095), .IN2(n6539), .IN3(\FIFO[93][0] ), .IN4(n6540), 
        .Q(n1555) );
  AO22X1 U1407 ( .IN1(n7078), .IN2(n6538), .IN3(\FIFO[93][1] ), .IN4(n6540), 
        .Q(n1556) );
  AO22X1 U1409 ( .IN1(n7056), .IN2(n6539), .IN3(\FIFO[93][3] ), .IN4(n6540), 
        .Q(n1558) );
  AO22X1 U1410 ( .IN1(n7045), .IN2(n6538), .IN3(\FIFO[93][4] ), .IN4(n6540), 
        .Q(n1559) );
  AO22X1 U1411 ( .IN1(n7034), .IN2(n6537), .IN3(\FIFO[93][5] ), .IN4(n6540), 
        .Q(n1560) );
  AO22X1 U1412 ( .IN1(n7023), .IN2(n6539), .IN3(\FIFO[93][6] ), .IN4(n6540), 
        .Q(n1561) );
  AO22X1 U1413 ( .IN1(n7012), .IN2(n6539), .IN3(\FIFO[93][7] ), .IN4(n6540), 
        .Q(n1562) );
  AO22X1 U1414 ( .IN1(n7001), .IN2(n6539), .IN3(\FIFO[93][8] ), .IN4(n6540), 
        .Q(n1563) );
  AO22X1 U1415 ( .IN1(n6990), .IN2(n6539), .IN3(\FIFO[93][9] ), .IN4(n6540), 
        .Q(n1564) );
  AO22X1 U1416 ( .IN1(n6979), .IN2(n6539), .IN3(\FIFO[93][10] ), .IN4(n6540), 
        .Q(n1565) );
  AO22X1 U1417 ( .IN1(n6968), .IN2(n6539), .IN3(\FIFO[93][11] ), .IN4(n6540), 
        .Q(n1566) );
  AO22X1 U1418 ( .IN1(n6957), .IN2(n6539), .IN3(\FIFO[93][12] ), .IN4(n6541), 
        .Q(n1567) );
  AO22X1 U1419 ( .IN1(n6946), .IN2(n6539), .IN3(\FIFO[93][13] ), .IN4(n6541), 
        .Q(n1568) );
  AO22X1 U1420 ( .IN1(n6935), .IN2(n6538), .IN3(\FIFO[93][14] ), .IN4(n6541), 
        .Q(n1569) );
  AO22X1 U1421 ( .IN1(n6924), .IN2(n6538), .IN3(\FIFO[93][15] ), .IN4(n6541), 
        .Q(n1570) );
  AO22X1 U1422 ( .IN1(n6913), .IN2(n6538), .IN3(\FIFO[93][16] ), .IN4(n6541), 
        .Q(n1571) );
  AO22X1 U1424 ( .IN1(n6891), .IN2(n6538), .IN3(\FIFO[93][18] ), .IN4(n6541), 
        .Q(n1573) );
  AO22X1 U1425 ( .IN1(n6880), .IN2(n6538), .IN3(\FIFO[93][19] ), .IN4(n6541), 
        .Q(n1574) );
  AO22X1 U1426 ( .IN1(n6869), .IN2(n6538), .IN3(\FIFO[93][20] ), .IN4(n6541), 
        .Q(n1575) );
  AO22X1 U1427 ( .IN1(n6858), .IN2(n6537), .IN3(\FIFO[93][21] ), .IN4(n6541), 
        .Q(n1576) );
  AO22X1 U1428 ( .IN1(n6847), .IN2(n6537), .IN3(\FIFO[93][22] ), .IN4(n6541), 
        .Q(n1577) );
  AO22X1 U1429 ( .IN1(n6836), .IN2(n6537), .IN3(\FIFO[93][23] ), .IN4(n6541), 
        .Q(n1578) );
  AO22X1 U1430 ( .IN1(n6825), .IN2(n6537), .IN3(\FIFO[93][24] ), .IN4(n6542), 
        .Q(n1579) );
  AO22X1 U1431 ( .IN1(n6814), .IN2(n6537), .IN3(\FIFO[93][25] ), .IN4(n6542), 
        .Q(n1580) );
  AO22X1 U1432 ( .IN1(n6803), .IN2(n6537), .IN3(\FIFO[93][26] ), .IN4(n6542), 
        .Q(n1581) );
  AO22X1 U1433 ( .IN1(n6792), .IN2(n6537), .IN3(\FIFO[93][27] ), .IN4(n6542), 
        .Q(n1582) );
  AO22X1 U1434 ( .IN1(n6781), .IN2(n6537), .IN3(\FIFO[93][28] ), .IN4(n6542), 
        .Q(n1583) );
  AO22X1 U1435 ( .IN1(n6770), .IN2(n6538), .IN3(\FIFO[93][29] ), .IN4(n6542), 
        .Q(n1584) );
  AO22X1 U1436 ( .IN1(n6759), .IN2(n6537), .IN3(\FIFO[93][30] ), .IN4(n6542), 
        .Q(n1585) );
  AO22X1 U1437 ( .IN1(n6748), .IN2(n6538), .IN3(\FIFO[93][31] ), .IN4(n6542), 
        .Q(n1586) );
  AO21X1 U1438 ( .IN1(n289), .IN2(n243), .IN3(n5975), .Q(n291) );
  AO22X1 U1439 ( .IN1(n7095), .IN2(n6533), .IN3(\FIFO[92][0] ), .IN4(n6534), 
        .Q(n1587) );
  AO22X1 U1440 ( .IN1(n7078), .IN2(n6533), .IN3(\FIFO[92][1] ), .IN4(n6534), 
        .Q(n1588) );
  AO22X1 U1441 ( .IN1(n7067), .IN2(n6533), .IN3(\FIFO[92][2] ), .IN4(n6534), 
        .Q(n1589) );
  AO22X1 U1442 ( .IN1(n7056), .IN2(n6533), .IN3(\FIFO[92][3] ), .IN4(n6534), 
        .Q(n1590) );
  AO22X1 U1443 ( .IN1(n7045), .IN2(n6533), .IN3(\FIFO[92][4] ), .IN4(n6534), 
        .Q(n1591) );
  AO22X1 U1444 ( .IN1(n7034), .IN2(n6533), .IN3(\FIFO[92][5] ), .IN4(n6534), 
        .Q(n1592) );
  AO22X1 U1445 ( .IN1(n7023), .IN2(n6533), .IN3(\FIFO[92][6] ), .IN4(n6534), 
        .Q(n1593) );
  AO22X1 U1446 ( .IN1(n7012), .IN2(n6532), .IN3(\FIFO[92][7] ), .IN4(n6534), 
        .Q(n1594) );
  AO22X1 U1447 ( .IN1(n7001), .IN2(n6532), .IN3(\FIFO[92][8] ), .IN4(n6534), 
        .Q(n1595) );
  AO22X1 U1448 ( .IN1(n6990), .IN2(n6532), .IN3(\FIFO[92][9] ), .IN4(n6534), 
        .Q(n1596) );
  AO22X1 U1449 ( .IN1(n6979), .IN2(n6532), .IN3(\FIFO[92][10] ), .IN4(n6534), 
        .Q(n1597) );
  AO22X1 U1450 ( .IN1(n6968), .IN2(n6532), .IN3(\FIFO[92][11] ), .IN4(n6534), 
        .Q(n1598) );
  AO22X1 U1451 ( .IN1(n6957), .IN2(n6532), .IN3(\FIFO[92][12] ), .IN4(n6535), 
        .Q(n1599) );
  AO22X1 U1452 ( .IN1(n6946), .IN2(n6532), .IN3(\FIFO[92][13] ), .IN4(n6535), 
        .Q(n1600) );
  AO22X1 U1453 ( .IN1(n6935), .IN2(n6531), .IN3(\FIFO[92][14] ), .IN4(n6535), 
        .Q(n1601) );
  AO22X1 U1454 ( .IN1(n6924), .IN2(n6531), .IN3(\FIFO[92][15] ), .IN4(n6535), 
        .Q(n1602) );
  AO22X1 U1455 ( .IN1(n6913), .IN2(n6531), .IN3(\FIFO[92][16] ), .IN4(n6535), 
        .Q(n1603) );
  AO22X1 U1456 ( .IN1(n6902), .IN2(n6531), .IN3(\FIFO[92][17] ), .IN4(n6535), 
        .Q(n1604) );
  AO22X1 U1457 ( .IN1(n6891), .IN2(n6531), .IN3(\FIFO[92][18] ), .IN4(n6535), 
        .Q(n1605) );
  AO22X1 U1458 ( .IN1(n6880), .IN2(n6531), .IN3(\FIFO[92][19] ), .IN4(n6535), 
        .Q(n1606) );
  AO22X1 U1459 ( .IN1(n6869), .IN2(n6531), .IN3(\FIFO[92][20] ), .IN4(n6535), 
        .Q(n1607) );
  AO22X1 U1460 ( .IN1(n6858), .IN2(n6533), .IN3(\FIFO[92][21] ), .IN4(n6535), 
        .Q(n1608) );
  AO22X1 U1461 ( .IN1(n6847), .IN2(n6532), .IN3(\FIFO[92][22] ), .IN4(n6535), 
        .Q(n1609) );
  AO22X1 U1462 ( .IN1(n6836), .IN2(n6531), .IN3(\FIFO[92][23] ), .IN4(n6535), 
        .Q(n1610) );
  AO22X1 U1463 ( .IN1(n6825), .IN2(n292), .IN3(\FIFO[92][24] ), .IN4(n6536), 
        .Q(n1611) );
  AO22X1 U1464 ( .IN1(n6814), .IN2(n292), .IN3(\FIFO[92][25] ), .IN4(n6536), 
        .Q(n1612) );
  AO22X1 U1465 ( .IN1(n6803), .IN2(n292), .IN3(\FIFO[92][26] ), .IN4(n6536), 
        .Q(n1613) );
  AO22X1 U1466 ( .IN1(n6792), .IN2(n6533), .IN3(\FIFO[92][27] ), .IN4(n6536), 
        .Q(n1614) );
  AO22X1 U1467 ( .IN1(n6781), .IN2(n6532), .IN3(\FIFO[92][28] ), .IN4(n6536), 
        .Q(n1615) );
  AO22X1 U1468 ( .IN1(n6770), .IN2(n6533), .IN3(\FIFO[92][29] ), .IN4(n6536), 
        .Q(n1616) );
  AO22X1 U1469 ( .IN1(n6759), .IN2(n6532), .IN3(\FIFO[92][30] ), .IN4(n6536), 
        .Q(n1617) );
  AO22X1 U1470 ( .IN1(n6748), .IN2(n6531), .IN3(\FIFO[92][31] ), .IN4(n6536), 
        .Q(n1618) );
  AO21X1 U1471 ( .IN1(n289), .IN2(n245), .IN3(n5974), .Q(n292) );
  AO22X1 U1496 ( .IN1(n6825), .IN2(n293), .IN3(\FIFO[91][24] ), .IN4(n6530), 
        .Q(n1643) );
  AO22X1 U1497 ( .IN1(n6814), .IN2(n293), .IN3(\FIFO[91][25] ), .IN4(n6530), 
        .Q(n1644) );
  AO22X1 U1498 ( .IN1(n6803), .IN2(n293), .IN3(\FIFO[91][26] ), .IN4(n6530), 
        .Q(n1645) );
  AO22X1 U1499 ( .IN1(n6792), .IN2(n6527), .IN3(\FIFO[91][27] ), .IN4(n6530), 
        .Q(n1646) );
  AO22X1 U1500 ( .IN1(n6781), .IN2(n6526), .IN3(\FIFO[91][28] ), .IN4(n6530), 
        .Q(n1647) );
  AO22X1 U1501 ( .IN1(n6770), .IN2(n6527), .IN3(\FIFO[91][29] ), .IN4(n6530), 
        .Q(n1648) );
  AO22X1 U1502 ( .IN1(n6759), .IN2(n6526), .IN3(\FIFO[91][30] ), .IN4(n6530), 
        .Q(n1649) );
  AO22X1 U1503 ( .IN1(n6748), .IN2(n6525), .IN3(\FIFO[91][31] ), .IN4(n6530), 
        .Q(n1650) );
  AO21X1 U1504 ( .IN1(n289), .IN2(n247), .IN3(flush), .Q(n293) );
  AO22X1 U1529 ( .IN1(n6825), .IN2(n294), .IN3(\FIFO[90][24] ), .IN4(n6524), 
        .Q(n1675) );
  AO22X1 U1530 ( .IN1(n6814), .IN2(n294), .IN3(\FIFO[90][25] ), .IN4(n6524), 
        .Q(n1676) );
  AO22X1 U1531 ( .IN1(n6803), .IN2(n294), .IN3(\FIFO[90][26] ), .IN4(n6524), 
        .Q(n1677) );
  AO22X1 U1532 ( .IN1(n6792), .IN2(n6521), .IN3(\FIFO[90][27] ), .IN4(n6524), 
        .Q(n1678) );
  AO22X1 U1533 ( .IN1(n6781), .IN2(n6521), .IN3(\FIFO[90][28] ), .IN4(n6524), 
        .Q(n1679) );
  AO22X1 U1534 ( .IN1(n6770), .IN2(n6520), .IN3(\FIFO[90][29] ), .IN4(n6524), 
        .Q(n1680) );
  AO22X1 U1535 ( .IN1(n6759), .IN2(n6519), .IN3(\FIFO[90][30] ), .IN4(n6524), 
        .Q(n1681) );
  AO22X1 U1536 ( .IN1(n6748), .IN2(n6520), .IN3(\FIFO[90][31] ), .IN4(n6524), 
        .Q(n1682) );
  AO21X1 U1537 ( .IN1(n289), .IN2(n249), .IN3(n5973), .Q(n294) );
  AO22X1 U1538 ( .IN1(n7095), .IN2(n6515), .IN3(\FIFO[89][0] ), .IN4(n6516), 
        .Q(n1683) );
  AO22X1 U1539 ( .IN1(n7078), .IN2(n6515), .IN3(\FIFO[89][1] ), .IN4(n6516), 
        .Q(n1684) );
  AO22X1 U1540 ( .IN1(n7067), .IN2(n6515), .IN3(\FIFO[89][2] ), .IN4(n6516), 
        .Q(n1685) );
  AO22X1 U1542 ( .IN1(n7045), .IN2(n6515), .IN3(\FIFO[89][4] ), .IN4(n6516), 
        .Q(n1687) );
  AO22X1 U1543 ( .IN1(n7034), .IN2(n6515), .IN3(\FIFO[89][5] ), .IN4(n6516), 
        .Q(n1688) );
  AO22X1 U1544 ( .IN1(n7023), .IN2(n6515), .IN3(\FIFO[89][6] ), .IN4(n6516), 
        .Q(n1689) );
  AO22X1 U1545 ( .IN1(n7012), .IN2(n6514), .IN3(\FIFO[89][7] ), .IN4(n6516), 
        .Q(n1690) );
  AO22X1 U1546 ( .IN1(n7001), .IN2(n6514), .IN3(\FIFO[89][8] ), .IN4(n6516), 
        .Q(n1691) );
  AO22X1 U1547 ( .IN1(n6990), .IN2(n6514), .IN3(\FIFO[89][9] ), .IN4(n6516), 
        .Q(n1692) );
  AO22X1 U1548 ( .IN1(n6979), .IN2(n6514), .IN3(\FIFO[89][10] ), .IN4(n6516), 
        .Q(n1693) );
  AO22X1 U1549 ( .IN1(n6968), .IN2(n6514), .IN3(\FIFO[89][11] ), .IN4(n6516), 
        .Q(n1694) );
  AO22X1 U1550 ( .IN1(n6957), .IN2(n6514), .IN3(\FIFO[89][12] ), .IN4(n6517), 
        .Q(n1695) );
  AO22X1 U1551 ( .IN1(n6946), .IN2(n6514), .IN3(\FIFO[89][13] ), .IN4(n6517), 
        .Q(n1696) );
  AO22X1 U1552 ( .IN1(n6935), .IN2(n6515), .IN3(\FIFO[89][14] ), .IN4(n6517), 
        .Q(n1697) );
  AO22X1 U1553 ( .IN1(n6924), .IN2(n6514), .IN3(\FIFO[89][15] ), .IN4(n6517), 
        .Q(n1698) );
  AO22X1 U1555 ( .IN1(n6902), .IN2(n6515), .IN3(\FIFO[89][17] ), .IN4(n6517), 
        .Q(n1700) );
  AO22X1 U1556 ( .IN1(n6891), .IN2(n6514), .IN3(\FIFO[89][18] ), .IN4(n6517), 
        .Q(n1701) );
  AO22X1 U1557 ( .IN1(n6880), .IN2(n6513), .IN3(\FIFO[89][19] ), .IN4(n6517), 
        .Q(n1702) );
  AO22X1 U1558 ( .IN1(n6869), .IN2(n6515), .IN3(\FIFO[89][20] ), .IN4(n6517), 
        .Q(n1703) );
  AO22X1 U1559 ( .IN1(n6858), .IN2(n6513), .IN3(\FIFO[89][21] ), .IN4(n6517), 
        .Q(n1704) );
  AO22X1 U1560 ( .IN1(n6847), .IN2(n6513), .IN3(\FIFO[89][22] ), .IN4(n6517), 
        .Q(n1705) );
  AO22X1 U1561 ( .IN1(n6836), .IN2(n6513), .IN3(\FIFO[89][23] ), .IN4(n6517), 
        .Q(n1706) );
  AO22X1 U1562 ( .IN1(n6825), .IN2(n6513), .IN3(\FIFO[89][24] ), .IN4(n6518), 
        .Q(n1707) );
  AO22X1 U1563 ( .IN1(n6814), .IN2(n6513), .IN3(\FIFO[89][25] ), .IN4(n6518), 
        .Q(n1708) );
  AO22X1 U1564 ( .IN1(n6803), .IN2(n6513), .IN3(\FIFO[89][26] ), .IN4(n6518), 
        .Q(n1709) );
  AO22X1 U1565 ( .IN1(n6792), .IN2(n6513), .IN3(\FIFO[89][27] ), .IN4(n6518), 
        .Q(n1710) );
  AO22X1 U1566 ( .IN1(n6781), .IN2(n6513), .IN3(\FIFO[89][28] ), .IN4(n6518), 
        .Q(n1711) );
  AO22X1 U1567 ( .IN1(n6770), .IN2(n6514), .IN3(\FIFO[89][29] ), .IN4(n6518), 
        .Q(n1712) );
  AO22X1 U1568 ( .IN1(n6759), .IN2(n6513), .IN3(\FIFO[89][30] ), .IN4(n6518), 
        .Q(n1713) );
  AO22X1 U1569 ( .IN1(n6748), .IN2(n6514), .IN3(\FIFO[89][31] ), .IN4(n6518), 
        .Q(n1714) );
  AO21X1 U1570 ( .IN1(n289), .IN2(n251), .IN3(n7359), .Q(n295) );
  AO22X1 U1571 ( .IN1(n7095), .IN2(n6509), .IN3(\FIFO[88][0] ), .IN4(n6510), 
        .Q(n1715) );
  AO22X1 U1572 ( .IN1(n7078), .IN2(n6508), .IN3(\FIFO[88][1] ), .IN4(n6510), 
        .Q(n1716) );
  AO22X1 U1573 ( .IN1(n7067), .IN2(n6507), .IN3(\FIFO[88][2] ), .IN4(n6510), 
        .Q(n1717) );
  AO22X1 U1574 ( .IN1(n7056), .IN2(n6509), .IN3(\FIFO[88][3] ), .IN4(n6510), 
        .Q(n1718) );
  AO22X1 U1576 ( .IN1(n7034), .IN2(n6507), .IN3(\FIFO[88][5] ), .IN4(n6510), 
        .Q(n1720) );
  AO22X1 U1577 ( .IN1(n7023), .IN2(n6509), .IN3(\FIFO[88][6] ), .IN4(n6510), 
        .Q(n1721) );
  AO22X1 U1578 ( .IN1(n7012), .IN2(n6509), .IN3(\FIFO[88][7] ), .IN4(n6510), 
        .Q(n1722) );
  AO22X1 U1579 ( .IN1(n7001), .IN2(n6509), .IN3(\FIFO[88][8] ), .IN4(n6510), 
        .Q(n1723) );
  AO22X1 U1580 ( .IN1(n6990), .IN2(n6509), .IN3(\FIFO[88][9] ), .IN4(n6510), 
        .Q(n1724) );
  AO22X1 U1581 ( .IN1(n6979), .IN2(n6509), .IN3(\FIFO[88][10] ), .IN4(n6510), 
        .Q(n1725) );
  AO22X1 U1582 ( .IN1(n6968), .IN2(n6509), .IN3(\FIFO[88][11] ), .IN4(n6510), 
        .Q(n1726) );
  AO22X1 U1583 ( .IN1(n6957), .IN2(n6509), .IN3(\FIFO[88][12] ), .IN4(n6511), 
        .Q(n1727) );
  AO22X1 U1584 ( .IN1(n6946), .IN2(n6509), .IN3(\FIFO[88][13] ), .IN4(n6511), 
        .Q(n1728) );
  AO22X1 U1585 ( .IN1(n6935), .IN2(n6508), .IN3(\FIFO[88][14] ), .IN4(n6511), 
        .Q(n1729) );
  AO22X1 U1586 ( .IN1(n6924), .IN2(n6508), .IN3(\FIFO[88][15] ), .IN4(n6511), 
        .Q(n1730) );
  AO22X1 U1587 ( .IN1(n6913), .IN2(n6508), .IN3(\FIFO[88][16] ), .IN4(n6511), 
        .Q(n1731) );
  AO22X1 U1588 ( .IN1(n6902), .IN2(n6508), .IN3(\FIFO[88][17] ), .IN4(n6511), 
        .Q(n1732) );
  AO22X1 U1589 ( .IN1(n6891), .IN2(n6508), .IN3(\FIFO[88][18] ), .IN4(n6511), 
        .Q(n1733) );
  AO22X1 U1590 ( .IN1(n6880), .IN2(n6508), .IN3(\FIFO[88][19] ), .IN4(n6511), 
        .Q(n1734) );
  AO22X1 U1591 ( .IN1(n6869), .IN2(n6508), .IN3(\FIFO[88][20] ), .IN4(n6511), 
        .Q(n1735) );
  AO22X1 U1592 ( .IN1(n6858), .IN2(n6507), .IN3(\FIFO[88][21] ), .IN4(n6511), 
        .Q(n1736) );
  AO22X1 U1593 ( .IN1(n6847), .IN2(n6507), .IN3(\FIFO[88][22] ), .IN4(n6511), 
        .Q(n1737) );
  AO22X1 U1594 ( .IN1(n6836), .IN2(n6507), .IN3(\FIFO[88][23] ), .IN4(n6511), 
        .Q(n1738) );
  AO22X1 U1595 ( .IN1(n6825), .IN2(n6507), .IN3(\FIFO[88][24] ), .IN4(n6512), 
        .Q(n1739) );
  AO22X1 U1596 ( .IN1(n6814), .IN2(n6507), .IN3(\FIFO[88][25] ), .IN4(n6512), 
        .Q(n1740) );
  AO22X1 U1597 ( .IN1(n6803), .IN2(n6507), .IN3(\FIFO[88][26] ), .IN4(n6512), 
        .Q(n1741) );
  AO22X1 U1598 ( .IN1(n6792), .IN2(n6507), .IN3(\FIFO[88][27] ), .IN4(n6512), 
        .Q(n1742) );
  AO22X1 U1599 ( .IN1(n6781), .IN2(n6507), .IN3(\FIFO[88][28] ), .IN4(n6512), 
        .Q(n1743) );
  AO22X1 U1600 ( .IN1(n6770), .IN2(n6508), .IN3(\FIFO[88][29] ), .IN4(n6512), 
        .Q(n1744) );
  AO22X1 U1601 ( .IN1(n6759), .IN2(n6507), .IN3(\FIFO[88][30] ), .IN4(n6512), 
        .Q(n1745) );
  AO22X1 U1602 ( .IN1(n6748), .IN2(n6508), .IN3(\FIFO[88][31] ), .IN4(n6512), 
        .Q(n1746) );
  AO21X1 U1603 ( .IN1(n289), .IN2(n253), .IN3(flush), .Q(n296) );
  AO22X1 U1628 ( .IN1(n6825), .IN2(n297), .IN3(\FIFO[87][24] ), .IN4(n6506), 
        .Q(n1771) );
  AO22X1 U1629 ( .IN1(n6814), .IN2(n297), .IN3(\FIFO[87][25] ), .IN4(n6506), 
        .Q(n1772) );
  AO22X1 U1630 ( .IN1(n6803), .IN2(n297), .IN3(\FIFO[87][26] ), .IN4(n6506), 
        .Q(n1773) );
  AO22X1 U1631 ( .IN1(n6792), .IN2(n6503), .IN3(\FIFO[87][27] ), .IN4(n6506), 
        .Q(n1774) );
  AO22X1 U1632 ( .IN1(n6781), .IN2(n6502), .IN3(\FIFO[87][28] ), .IN4(n6506), 
        .Q(n1775) );
  AO22X1 U1633 ( .IN1(n6770), .IN2(n6503), .IN3(\FIFO[87][29] ), .IN4(n6506), 
        .Q(n1776) );
  AO22X1 U1634 ( .IN1(n6759), .IN2(n6502), .IN3(\FIFO[87][30] ), .IN4(n6506), 
        .Q(n1777) );
  AO22X1 U1635 ( .IN1(n6748), .IN2(n6501), .IN3(\FIFO[87][31] ), .IN4(n6506), 
        .Q(n1778) );
  AO21X1 U1636 ( .IN1(n289), .IN2(n255), .IN3(n5973), .Q(n297) );
  AO22X1 U1661 ( .IN1(n6825), .IN2(n298), .IN3(\FIFO[86][24] ), .IN4(n6500), 
        .Q(n1803) );
  AO22X1 U1662 ( .IN1(n6814), .IN2(n298), .IN3(\FIFO[86][25] ), .IN4(n6500), 
        .Q(n1804) );
  AO22X1 U1663 ( .IN1(n6803), .IN2(n298), .IN3(\FIFO[86][26] ), .IN4(n6500), 
        .Q(n1805) );
  AO22X1 U1664 ( .IN1(n6792), .IN2(n6497), .IN3(\FIFO[86][27] ), .IN4(n6500), 
        .Q(n1806) );
  AO22X1 U1665 ( .IN1(n6781), .IN2(n6496), .IN3(\FIFO[86][28] ), .IN4(n6500), 
        .Q(n1807) );
  AO22X1 U1666 ( .IN1(n6770), .IN2(n6497), .IN3(\FIFO[86][29] ), .IN4(n6500), 
        .Q(n1808) );
  AO22X1 U1667 ( .IN1(n6759), .IN2(n6496), .IN3(\FIFO[86][30] ), .IN4(n6500), 
        .Q(n1809) );
  AO22X1 U1668 ( .IN1(n6748), .IN2(n6495), .IN3(\FIFO[86][31] ), .IN4(n6500), 
        .Q(n1810) );
  AO21X1 U1669 ( .IN1(n289), .IN2(n257), .IN3(n7359), .Q(n298) );
  AO22X1 U1670 ( .IN1(n7095), .IN2(n6491), .IN3(\FIFO[85][0] ), .IN4(n6492), 
        .Q(n1811) );
  AO22X1 U1671 ( .IN1(n7078), .IN2(n6491), .IN3(\FIFO[85][1] ), .IN4(n6492), 
        .Q(n1812) );
  AO22X1 U1672 ( .IN1(n7067), .IN2(n6491), .IN3(\FIFO[85][2] ), .IN4(n6492), 
        .Q(n1813) );
  AO22X1 U1673 ( .IN1(n7056), .IN2(n6491), .IN3(\FIFO[85][3] ), .IN4(n6492), 
        .Q(n1814) );
  AO22X1 U1674 ( .IN1(n7045), .IN2(n6491), .IN3(\FIFO[85][4] ), .IN4(n6492), 
        .Q(n1815) );
  AO22X1 U1675 ( .IN1(n7034), .IN2(n6491), .IN3(\FIFO[85][5] ), .IN4(n6492), 
        .Q(n1816) );
  AO22X1 U1676 ( .IN1(n7023), .IN2(n6491), .IN3(\FIFO[85][6] ), .IN4(n6492), 
        .Q(n1817) );
  AO22X1 U1677 ( .IN1(n7012), .IN2(n6490), .IN3(\FIFO[85][7] ), .IN4(n6492), 
        .Q(n1818) );
  AO22X1 U1678 ( .IN1(n7001), .IN2(n6490), .IN3(\FIFO[85][8] ), .IN4(n6492), 
        .Q(n1819) );
  AO22X1 U1679 ( .IN1(n6990), .IN2(n6490), .IN3(\FIFO[85][9] ), .IN4(n6492), 
        .Q(n1820) );
  AO22X1 U1680 ( .IN1(n6979), .IN2(n6490), .IN3(\FIFO[85][10] ), .IN4(n6492), 
        .Q(n1821) );
  AO22X1 U1681 ( .IN1(n6968), .IN2(n6490), .IN3(\FIFO[85][11] ), .IN4(n6492), 
        .Q(n1822) );
  AO22X1 U1682 ( .IN1(n6957), .IN2(n6490), .IN3(\FIFO[85][12] ), .IN4(n6493), 
        .Q(n1823) );
  AO22X1 U1683 ( .IN1(n6946), .IN2(n6490), .IN3(\FIFO[85][13] ), .IN4(n6493), 
        .Q(n1824) );
  AO22X1 U1684 ( .IN1(n6935), .IN2(n6489), .IN3(\FIFO[85][14] ), .IN4(n6493), 
        .Q(n1825) );
  AO22X1 U1685 ( .IN1(n6924), .IN2(n6489), .IN3(\FIFO[85][15] ), .IN4(n6493), 
        .Q(n1826) );
  AO22X1 U1686 ( .IN1(n6913), .IN2(n6489), .IN3(\FIFO[85][16] ), .IN4(n6493), 
        .Q(n1827) );
  AO22X1 U1687 ( .IN1(n6902), .IN2(n6489), .IN3(\FIFO[85][17] ), .IN4(n6493), 
        .Q(n1828) );
  AO22X1 U1688 ( .IN1(n6891), .IN2(n6489), .IN3(\FIFO[85][18] ), .IN4(n6493), 
        .Q(n1829) );
  AO22X1 U1689 ( .IN1(n6880), .IN2(n6489), .IN3(\FIFO[85][19] ), .IN4(n6493), 
        .Q(n1830) );
  AO22X1 U1690 ( .IN1(n6869), .IN2(n6489), .IN3(\FIFO[85][20] ), .IN4(n6493), 
        .Q(n1831) );
  AO22X1 U1691 ( .IN1(n6858), .IN2(n6491), .IN3(\FIFO[85][21] ), .IN4(n6493), 
        .Q(n1832) );
  AO22X1 U1692 ( .IN1(n6847), .IN2(n6490), .IN3(\FIFO[85][22] ), .IN4(n6493), 
        .Q(n1833) );
  AO22X1 U1693 ( .IN1(n6836), .IN2(n6489), .IN3(\FIFO[85][23] ), .IN4(n6493), 
        .Q(n1834) );
  AO22X1 U1694 ( .IN1(n6825), .IN2(n299), .IN3(\FIFO[85][24] ), .IN4(n6494), 
        .Q(n1835) );
  AO22X1 U1695 ( .IN1(n6814), .IN2(n299), .IN3(\FIFO[85][25] ), .IN4(n6494), 
        .Q(n1836) );
  AO22X1 U1696 ( .IN1(n6803), .IN2(n299), .IN3(\FIFO[85][26] ), .IN4(n6494), 
        .Q(n1837) );
  AO22X1 U1697 ( .IN1(n6792), .IN2(n6491), .IN3(\FIFO[85][27] ), .IN4(n6494), 
        .Q(n1838) );
  AO22X1 U1698 ( .IN1(n6781), .IN2(n6491), .IN3(\FIFO[85][28] ), .IN4(n6494), 
        .Q(n1839) );
  AO22X1 U1699 ( .IN1(n6770), .IN2(n6490), .IN3(\FIFO[85][29] ), .IN4(n6494), 
        .Q(n1840) );
  AO22X1 U1700 ( .IN1(n6759), .IN2(n6489), .IN3(\FIFO[85][30] ), .IN4(n6494), 
        .Q(n1841) );
  AO22X1 U1701 ( .IN1(n6748), .IN2(n6490), .IN3(\FIFO[85][31] ), .IN4(n6494), 
        .Q(n1842) );
  AO21X1 U1702 ( .IN1(n289), .IN2(n259), .IN3(flush), .Q(n299) );
  AO22X1 U1703 ( .IN1(n7095), .IN2(n6485), .IN3(\FIFO[84][0] ), .IN4(n6486), 
        .Q(n1843) );
  AO22X1 U1704 ( .IN1(n7078), .IN2(n6485), .IN3(\FIFO[84][1] ), .IN4(n6486), 
        .Q(n1844) );
  AO22X1 U1705 ( .IN1(n7067), .IN2(n6485), .IN3(\FIFO[84][2] ), .IN4(n6486), 
        .Q(n1845) );
  AO22X1 U1706 ( .IN1(n7056), .IN2(n6485), .IN3(\FIFO[84][3] ), .IN4(n6486), 
        .Q(n1846) );
  AO22X1 U1707 ( .IN1(n7045), .IN2(n6485), .IN3(\FIFO[84][4] ), .IN4(n6486), 
        .Q(n1847) );
  AO22X1 U1709 ( .IN1(n7023), .IN2(n6485), .IN3(\FIFO[84][6] ), .IN4(n6486), 
        .Q(n1849) );
  AO22X1 U1710 ( .IN1(n7012), .IN2(n6484), .IN3(\FIFO[84][7] ), .IN4(n6486), 
        .Q(n1850) );
  AO22X1 U1711 ( .IN1(n7001), .IN2(n6484), .IN3(\FIFO[84][8] ), .IN4(n6486), 
        .Q(n1851) );
  AO22X1 U1712 ( .IN1(n6990), .IN2(n6484), .IN3(\FIFO[84][9] ), .IN4(n6486), 
        .Q(n1852) );
  AO22X1 U1713 ( .IN1(n6979), .IN2(n6484), .IN3(\FIFO[84][10] ), .IN4(n6486), 
        .Q(n1853) );
  AO22X1 U1714 ( .IN1(n6968), .IN2(n6484), .IN3(\FIFO[84][11] ), .IN4(n6486), 
        .Q(n1854) );
  AO22X1 U1715 ( .IN1(n6957), .IN2(n6484), .IN3(\FIFO[84][12] ), .IN4(n6487), 
        .Q(n1855) );
  AO22X1 U1716 ( .IN1(n6946), .IN2(n6484), .IN3(\FIFO[84][13] ), .IN4(n6487), 
        .Q(n1856) );
  AO22X1 U1717 ( .IN1(n6935), .IN2(n6485), .IN3(\FIFO[84][14] ), .IN4(n6487), 
        .Q(n1857) );
  AO22X1 U1718 ( .IN1(n6924), .IN2(n6484), .IN3(\FIFO[84][15] ), .IN4(n6487), 
        .Q(n1858) );
  AO22X1 U1719 ( .IN1(n6913), .IN2(n6483), .IN3(\FIFO[84][16] ), .IN4(n6487), 
        .Q(n1859) );
  AO22X1 U1720 ( .IN1(n6902), .IN2(n6485), .IN3(\FIFO[84][17] ), .IN4(n6487), 
        .Q(n1860) );
  AO22X1 U1722 ( .IN1(n6880), .IN2(n6483), .IN3(\FIFO[84][19] ), .IN4(n6487), 
        .Q(n1862) );
  AO22X1 U1723 ( .IN1(n6869), .IN2(n6485), .IN3(\FIFO[84][20] ), .IN4(n6487), 
        .Q(n1863) );
  AO22X1 U1724 ( .IN1(n6858), .IN2(n6483), .IN3(\FIFO[84][21] ), .IN4(n6487), 
        .Q(n1864) );
  AO22X1 U1725 ( .IN1(n6847), .IN2(n6483), .IN3(\FIFO[84][22] ), .IN4(n6487), 
        .Q(n1865) );
  AO22X1 U1726 ( .IN1(n6836), .IN2(n6483), .IN3(\FIFO[84][23] ), .IN4(n6487), 
        .Q(n1866) );
  AO22X1 U1727 ( .IN1(n6825), .IN2(n6483), .IN3(\FIFO[84][24] ), .IN4(n6488), 
        .Q(n1867) );
  AO22X1 U1728 ( .IN1(n6814), .IN2(n6483), .IN3(\FIFO[84][25] ), .IN4(n6488), 
        .Q(n1868) );
  AO22X1 U1729 ( .IN1(n6803), .IN2(n6483), .IN3(\FIFO[84][26] ), .IN4(n6488), 
        .Q(n1869) );
  AO22X1 U1730 ( .IN1(n6792), .IN2(n6483), .IN3(\FIFO[84][27] ), .IN4(n6488), 
        .Q(n1870) );
  AO22X1 U1731 ( .IN1(n6781), .IN2(n6483), .IN3(\FIFO[84][28] ), .IN4(n6488), 
        .Q(n1871) );
  AO22X1 U1732 ( .IN1(n6770), .IN2(n6484), .IN3(\FIFO[84][29] ), .IN4(n6488), 
        .Q(n1872) );
  AO22X1 U1733 ( .IN1(n6759), .IN2(n6483), .IN3(\FIFO[84][30] ), .IN4(n6488), 
        .Q(n1873) );
  AO22X1 U1734 ( .IN1(n6748), .IN2(n6484), .IN3(\FIFO[84][31] ), .IN4(n6488), 
        .Q(n1874) );
  AO21X1 U1735 ( .IN1(n289), .IN2(n261), .IN3(n5973), .Q(n300) );
  AO22X1 U1760 ( .IN1(n6824), .IN2(n6477), .IN3(\FIFO[83][24] ), .IN4(n6482), 
        .Q(n1899) );
  AO22X1 U1761 ( .IN1(n6813), .IN2(n6477), .IN3(\FIFO[83][25] ), .IN4(n6482), 
        .Q(n1900) );
  AO22X1 U1762 ( .IN1(n6802), .IN2(n6477), .IN3(\FIFO[83][26] ), .IN4(n6482), 
        .Q(n1901) );
  AO22X1 U1763 ( .IN1(n6791), .IN2(n6477), .IN3(\FIFO[83][27] ), .IN4(n6482), 
        .Q(n1902) );
  AO22X1 U1764 ( .IN1(n6780), .IN2(n6477), .IN3(\FIFO[83][28] ), .IN4(n6482), 
        .Q(n1903) );
  AO22X1 U1765 ( .IN1(n6769), .IN2(n6478), .IN3(\FIFO[83][29] ), .IN4(n6482), 
        .Q(n1904) );
  AO22X1 U1766 ( .IN1(n6758), .IN2(n6477), .IN3(\FIFO[83][30] ), .IN4(n6482), 
        .Q(n1905) );
  AO22X1 U1767 ( .IN1(n6747), .IN2(n6478), .IN3(\FIFO[83][31] ), .IN4(n6482), 
        .Q(n1906) );
  AO21X1 U1768 ( .IN1(n289), .IN2(n263), .IN3(n7359), .Q(n301) );
  AO22X1 U1793 ( .IN1(n6824), .IN2(n302), .IN3(\FIFO[82][24] ), .IN4(n6476), 
        .Q(n1931) );
  AO22X1 U1794 ( .IN1(n6813), .IN2(n302), .IN3(\FIFO[82][25] ), .IN4(n6476), 
        .Q(n1932) );
  AO22X1 U1795 ( .IN1(n6802), .IN2(n302), .IN3(\FIFO[82][26] ), .IN4(n6476), 
        .Q(n1933) );
  AO22X1 U1796 ( .IN1(n6791), .IN2(n6473), .IN3(\FIFO[82][27] ), .IN4(n6476), 
        .Q(n1934) );
  AO22X1 U1797 ( .IN1(n6780), .IN2(n6472), .IN3(\FIFO[82][28] ), .IN4(n6476), 
        .Q(n1935) );
  AO22X1 U1798 ( .IN1(n6769), .IN2(n6473), .IN3(\FIFO[82][29] ), .IN4(n6476), 
        .Q(n1936) );
  AO22X1 U1799 ( .IN1(n6758), .IN2(n6472), .IN3(\FIFO[82][30] ), .IN4(n6476), 
        .Q(n1937) );
  AO22X1 U1800 ( .IN1(n6747), .IN2(n6471), .IN3(\FIFO[82][31] ), .IN4(n6476), 
        .Q(n1938) );
  AO21X1 U1801 ( .IN1(n289), .IN2(n265), .IN3(flush), .Q(n302) );
  AO22X1 U1802 ( .IN1(n7094), .IN2(n6467), .IN3(\FIFO[81][0] ), .IN4(n6468), 
        .Q(n1939) );
  AO22X1 U1803 ( .IN1(n7077), .IN2(n6467), .IN3(\FIFO[81][1] ), .IN4(n6468), 
        .Q(n1940) );
  AO22X1 U1804 ( .IN1(n7066), .IN2(n6467), .IN3(\FIFO[81][2] ), .IN4(n6468), 
        .Q(n1941) );
  AO22X1 U1805 ( .IN1(n7055), .IN2(n6467), .IN3(\FIFO[81][3] ), .IN4(n6468), 
        .Q(n1942) );
  AO22X1 U1806 ( .IN1(n7044), .IN2(n6467), .IN3(\FIFO[81][4] ), .IN4(n6468), 
        .Q(n1943) );
  AO22X1 U1807 ( .IN1(n7033), .IN2(n6467), .IN3(\FIFO[81][5] ), .IN4(n6468), 
        .Q(n1944) );
  AO22X1 U1808 ( .IN1(n7022), .IN2(n6467), .IN3(\FIFO[81][6] ), .IN4(n6468), 
        .Q(n1945) );
  AO22X1 U1809 ( .IN1(n7011), .IN2(n6466), .IN3(\FIFO[81][7] ), .IN4(n6468), 
        .Q(n1946) );
  AO22X1 U1810 ( .IN1(n7000), .IN2(n6466), .IN3(\FIFO[81][8] ), .IN4(n6468), 
        .Q(n1947) );
  AO22X1 U1811 ( .IN1(n6989), .IN2(n6466), .IN3(\FIFO[81][9] ), .IN4(n6468), 
        .Q(n1948) );
  AO22X1 U1812 ( .IN1(n6978), .IN2(n6466), .IN3(\FIFO[81][10] ), .IN4(n6468), 
        .Q(n1949) );
  AO22X1 U1813 ( .IN1(n6967), .IN2(n6466), .IN3(\FIFO[81][11] ), .IN4(n6468), 
        .Q(n1950) );
  AO22X1 U1814 ( .IN1(n6956), .IN2(n6466), .IN3(\FIFO[81][12] ), .IN4(n6469), 
        .Q(n1951) );
  AO22X1 U1815 ( .IN1(n6945), .IN2(n6466), .IN3(\FIFO[81][13] ), .IN4(n6469), 
        .Q(n1952) );
  AO22X1 U1816 ( .IN1(n6934), .IN2(n6465), .IN3(\FIFO[81][14] ), .IN4(n6469), 
        .Q(n1953) );
  AO22X1 U1817 ( .IN1(n6923), .IN2(n6465), .IN3(\FIFO[81][15] ), .IN4(n6469), 
        .Q(n1954) );
  AO22X1 U1818 ( .IN1(n6912), .IN2(n6465), .IN3(\FIFO[81][16] ), .IN4(n6469), 
        .Q(n1955) );
  AO22X1 U1819 ( .IN1(n6901), .IN2(n6465), .IN3(\FIFO[81][17] ), .IN4(n6469), 
        .Q(n1956) );
  AO22X1 U1820 ( .IN1(n6890), .IN2(n6465), .IN3(\FIFO[81][18] ), .IN4(n6469), 
        .Q(n1957) );
  AO22X1 U1821 ( .IN1(n6879), .IN2(n6465), .IN3(\FIFO[81][19] ), .IN4(n6469), 
        .Q(n1958) );
  AO22X1 U1822 ( .IN1(n6868), .IN2(n6465), .IN3(\FIFO[81][20] ), .IN4(n6469), 
        .Q(n1959) );
  AO22X1 U1823 ( .IN1(n6857), .IN2(n6467), .IN3(\FIFO[81][21] ), .IN4(n6469), 
        .Q(n1960) );
  AO22X1 U1824 ( .IN1(n6846), .IN2(n6466), .IN3(\FIFO[81][22] ), .IN4(n6469), 
        .Q(n1961) );
  AO22X1 U1825 ( .IN1(n6835), .IN2(n6465), .IN3(\FIFO[81][23] ), .IN4(n6469), 
        .Q(n1962) );
  AO22X1 U1826 ( .IN1(n6824), .IN2(n303), .IN3(\FIFO[81][24] ), .IN4(n6470), 
        .Q(n1963) );
  AO22X1 U1827 ( .IN1(n6813), .IN2(n303), .IN3(\FIFO[81][25] ), .IN4(n6470), 
        .Q(n1964) );
  AO22X1 U1828 ( .IN1(n6802), .IN2(n303), .IN3(\FIFO[81][26] ), .IN4(n6470), 
        .Q(n1965) );
  AO22X1 U1829 ( .IN1(n6791), .IN2(n6467), .IN3(\FIFO[81][27] ), .IN4(n6470), 
        .Q(n1966) );
  AO22X1 U1830 ( .IN1(n6780), .IN2(n6466), .IN3(\FIFO[81][28] ), .IN4(n6470), 
        .Q(n1967) );
  AO22X1 U1831 ( .IN1(n6769), .IN2(n6467), .IN3(\FIFO[81][29] ), .IN4(n6470), 
        .Q(n1968) );
  AO22X1 U1832 ( .IN1(n6758), .IN2(n6466), .IN3(\FIFO[81][30] ), .IN4(n6470), 
        .Q(n1969) );
  AO22X1 U1833 ( .IN1(n6747), .IN2(n6465), .IN3(\FIFO[81][31] ), .IN4(n6470), 
        .Q(n1970) );
  AO21X1 U1834 ( .IN1(n289), .IN2(n267), .IN3(n5973), .Q(n303) );
  AO22X1 U1835 ( .IN1(n7094), .IN2(n6461), .IN3(\FIFO[80][0] ), .IN4(n6462), 
        .Q(n1971) );
  AO22X1 U1836 ( .IN1(n7077), .IN2(n6461), .IN3(\FIFO[80][1] ), .IN4(n6462), 
        .Q(n1972) );
  AO22X1 U1837 ( .IN1(n7066), .IN2(n6461), .IN3(\FIFO[80][2] ), .IN4(n6462), 
        .Q(n1973) );
  AO22X1 U1838 ( .IN1(n7055), .IN2(n6461), .IN3(\FIFO[80][3] ), .IN4(n6462), 
        .Q(n1974) );
  AO22X1 U1839 ( .IN1(n7044), .IN2(n6461), .IN3(\FIFO[80][4] ), .IN4(n6462), 
        .Q(n1975) );
  AO22X1 U1840 ( .IN1(n7033), .IN2(n6461), .IN3(\FIFO[80][5] ), .IN4(n6462), 
        .Q(n1976) );
  AO22X1 U1841 ( .IN1(n7022), .IN2(n6461), .IN3(\FIFO[80][6] ), .IN4(n6462), 
        .Q(n1977) );
  AO22X1 U1842 ( .IN1(n7011), .IN2(n6460), .IN3(\FIFO[80][7] ), .IN4(n6462), 
        .Q(n1978) );
  AO22X1 U1843 ( .IN1(n7000), .IN2(n6460), .IN3(\FIFO[80][8] ), .IN4(n6462), 
        .Q(n1979) );
  AO22X1 U1844 ( .IN1(n6989), .IN2(n6460), .IN3(\FIFO[80][9] ), .IN4(n6462), 
        .Q(n1980) );
  AO22X1 U1845 ( .IN1(n6978), .IN2(n6460), .IN3(\FIFO[80][10] ), .IN4(n6462), 
        .Q(n1981) );
  AO22X1 U1846 ( .IN1(n6967), .IN2(n6460), .IN3(\FIFO[80][11] ), .IN4(n6462), 
        .Q(n1982) );
  AO22X1 U1847 ( .IN1(n6956), .IN2(n6460), .IN3(\FIFO[80][12] ), .IN4(n6463), 
        .Q(n1983) );
  AO22X1 U1848 ( .IN1(n6945), .IN2(n6460), .IN3(\FIFO[80][13] ), .IN4(n6463), 
        .Q(n1984) );
  AO22X1 U1849 ( .IN1(n6934), .IN2(n6459), .IN3(\FIFO[80][14] ), .IN4(n6463), 
        .Q(n1985) );
  AO22X1 U1850 ( .IN1(n6923), .IN2(n6459), .IN3(\FIFO[80][15] ), .IN4(n6463), 
        .Q(n1986) );
  AO22X1 U1851 ( .IN1(n6912), .IN2(n6459), .IN3(\FIFO[80][16] ), .IN4(n6463), 
        .Q(n1987) );
  AO22X1 U1852 ( .IN1(n6901), .IN2(n6459), .IN3(\FIFO[80][17] ), .IN4(n6463), 
        .Q(n1988) );
  AO22X1 U1853 ( .IN1(n6890), .IN2(n6459), .IN3(\FIFO[80][18] ), .IN4(n6463), 
        .Q(n1989) );
  AO22X1 U1854 ( .IN1(n6879), .IN2(n6459), .IN3(\FIFO[80][19] ), .IN4(n6463), 
        .Q(n1990) );
  AO22X1 U1855 ( .IN1(n6868), .IN2(n6459), .IN3(\FIFO[80][20] ), .IN4(n6463), 
        .Q(n1991) );
  AO22X1 U1856 ( .IN1(n6857), .IN2(n6461), .IN3(\FIFO[80][21] ), .IN4(n6463), 
        .Q(n1992) );
  AO22X1 U1857 ( .IN1(n6846), .IN2(n6460), .IN3(\FIFO[80][22] ), .IN4(n6463), 
        .Q(n1993) );
  AO22X1 U1858 ( .IN1(n6835), .IN2(n6459), .IN3(\FIFO[80][23] ), .IN4(n6463), 
        .Q(n1994) );
  AO22X1 U1859 ( .IN1(n6824), .IN2(n304), .IN3(\FIFO[80][24] ), .IN4(n6464), 
        .Q(n1995) );
  AO22X1 U1860 ( .IN1(n6813), .IN2(n304), .IN3(\FIFO[80][25] ), .IN4(n6464), 
        .Q(n1996) );
  AO22X1 U1861 ( .IN1(n6802), .IN2(n304), .IN3(\FIFO[80][26] ), .IN4(n6464), 
        .Q(n1997) );
  AO22X1 U1862 ( .IN1(n6791), .IN2(n6461), .IN3(\FIFO[80][27] ), .IN4(n6464), 
        .Q(n1998) );
  AO22X1 U1863 ( .IN1(n6780), .IN2(n6461), .IN3(\FIFO[80][28] ), .IN4(n6464), 
        .Q(n1999) );
  AO22X1 U1864 ( .IN1(n6769), .IN2(n6460), .IN3(\FIFO[80][29] ), .IN4(n6464), 
        .Q(n2000) );
  AO22X1 U1865 ( .IN1(n6758), .IN2(n6459), .IN3(\FIFO[80][30] ), .IN4(n6464), 
        .Q(n2001) );
  AO22X1 U1866 ( .IN1(n6747), .IN2(n6460), .IN3(\FIFO[80][31] ), .IN4(n6464), 
        .Q(n2002) );
  AO21X1 U1867 ( .IN1(n289), .IN2(n269), .IN3(n7359), .Q(n304) );
  AO22X1 U1893 ( .IN1(n6824), .IN2(n305), .IN3(\FIFO[79][24] ), .IN4(n6458), 
        .Q(n2027) );
  AO22X1 U1894 ( .IN1(n6813), .IN2(n305), .IN3(\FIFO[79][25] ), .IN4(n6458), 
        .Q(n2028) );
  AO22X1 U1895 ( .IN1(n6802), .IN2(n305), .IN3(\FIFO[79][26] ), .IN4(n6458), 
        .Q(n2029) );
  AO22X1 U1896 ( .IN1(n6791), .IN2(n6455), .IN3(\FIFO[79][27] ), .IN4(n6458), 
        .Q(n2030) );
  AO22X1 U1897 ( .IN1(n6780), .IN2(n6454), .IN3(\FIFO[79][28] ), .IN4(n6458), 
        .Q(n2031) );
  AO22X1 U1898 ( .IN1(n6769), .IN2(n6455), .IN3(\FIFO[79][29] ), .IN4(n6458), 
        .Q(n2032) );
  AO22X1 U1899 ( .IN1(n6758), .IN2(n6454), .IN3(\FIFO[79][30] ), .IN4(n6458), 
        .Q(n2033) );
  AO22X1 U1900 ( .IN1(n6747), .IN2(n6453), .IN3(\FIFO[79][31] ), .IN4(n6458), 
        .Q(n2034) );
  AO21X1 U1901 ( .IN1(n306), .IN2(n238), .IN3(flush), .Q(n305) );
  AO22X1 U1926 ( .IN1(n6824), .IN2(n307), .IN3(\FIFO[78][24] ), .IN4(n6452), 
        .Q(n2059) );
  AO22X1 U1927 ( .IN1(n6813), .IN2(n307), .IN3(\FIFO[78][25] ), .IN4(n6452), 
        .Q(n2060) );
  AO22X1 U1928 ( .IN1(n6802), .IN2(n307), .IN3(\FIFO[78][26] ), .IN4(n6452), 
        .Q(n2061) );
  AO22X1 U1929 ( .IN1(n6791), .IN2(n6449), .IN3(\FIFO[78][27] ), .IN4(n6452), 
        .Q(n2062) );
  AO22X1 U1930 ( .IN1(n6780), .IN2(n6449), .IN3(\FIFO[78][28] ), .IN4(n6452), 
        .Q(n2063) );
  AO22X1 U1931 ( .IN1(n6769), .IN2(n6448), .IN3(\FIFO[78][29] ), .IN4(n6452), 
        .Q(n2064) );
  AO22X1 U1932 ( .IN1(n6758), .IN2(n6447), .IN3(\FIFO[78][30] ), .IN4(n6452), 
        .Q(n2065) );
  AO22X1 U1933 ( .IN1(n6747), .IN2(n6448), .IN3(\FIFO[78][31] ), .IN4(n6452), 
        .Q(n2066) );
  AO21X1 U1934 ( .IN1(n306), .IN2(n241), .IN3(n5973), .Q(n307) );
  AO22X1 U1935 ( .IN1(n7094), .IN2(n6443), .IN3(\FIFO[77][0] ), .IN4(n6444), 
        .Q(n2067) );
  AO22X1 U1936 ( .IN1(n7077), .IN2(n6443), .IN3(\FIFO[77][1] ), .IN4(n6444), 
        .Q(n2068) );
  AO22X1 U1937 ( .IN1(n7066), .IN2(n6443), .IN3(\FIFO[77][2] ), .IN4(n6444), 
        .Q(n2069) );
  AO22X1 U1938 ( .IN1(n7055), .IN2(n6443), .IN3(\FIFO[77][3] ), .IN4(n6444), 
        .Q(n2070) );
  AO22X1 U1939 ( .IN1(n7044), .IN2(n6443), .IN3(\FIFO[77][4] ), .IN4(n6444), 
        .Q(n2071) );
  AO22X1 U1940 ( .IN1(n7033), .IN2(n6443), .IN3(\FIFO[77][5] ), .IN4(n6444), 
        .Q(n2072) );
  AO22X1 U1941 ( .IN1(n7022), .IN2(n6443), .IN3(\FIFO[77][6] ), .IN4(n6444), 
        .Q(n2073) );
  AO22X1 U1943 ( .IN1(n7000), .IN2(n6442), .IN3(\FIFO[77][8] ), .IN4(n6444), 
        .Q(n2075) );
  AO22X1 U1944 ( .IN1(n6989), .IN2(n6442), .IN3(\FIFO[77][9] ), .IN4(n6444), 
        .Q(n2076) );
  AO22X1 U1945 ( .IN1(n6978), .IN2(n6442), .IN3(\FIFO[77][10] ), .IN4(n6444), 
        .Q(n2077) );
  AO22X1 U1946 ( .IN1(n6967), .IN2(n6442), .IN3(\FIFO[77][11] ), .IN4(n6444), 
        .Q(n2078) );
  AO22X1 U1947 ( .IN1(n6956), .IN2(n6442), .IN3(\FIFO[77][12] ), .IN4(n6445), 
        .Q(n2079) );
  AO22X1 U1948 ( .IN1(n6945), .IN2(n6442), .IN3(\FIFO[77][13] ), .IN4(n6445), 
        .Q(n2080) );
  AO22X1 U1949 ( .IN1(n6934), .IN2(n6443), .IN3(\FIFO[77][14] ), .IN4(n6445), 
        .Q(n2081) );
  AO22X1 U1950 ( .IN1(n6923), .IN2(n6442), .IN3(\FIFO[77][15] ), .IN4(n6445), 
        .Q(n2082) );
  AO22X1 U1951 ( .IN1(n6912), .IN2(n6441), .IN3(\FIFO[77][16] ), .IN4(n6445), 
        .Q(n2083) );
  AO22X1 U1952 ( .IN1(n6901), .IN2(n6443), .IN3(\FIFO[77][17] ), .IN4(n6445), 
        .Q(n2084) );
  AO22X1 U1953 ( .IN1(n6890), .IN2(n6442), .IN3(\FIFO[77][18] ), .IN4(n6445), 
        .Q(n2085) );
  AO22X1 U1955 ( .IN1(n6868), .IN2(n6443), .IN3(\FIFO[77][20] ), .IN4(n6445), 
        .Q(n2087) );
  AO22X1 U1956 ( .IN1(n6857), .IN2(n6441), .IN3(\FIFO[77][21] ), .IN4(n6445), 
        .Q(n2088) );
  AO22X1 U1957 ( .IN1(n6846), .IN2(n6441), .IN3(\FIFO[77][22] ), .IN4(n6445), 
        .Q(n2089) );
  AO22X1 U1958 ( .IN1(n6835), .IN2(n6441), .IN3(\FIFO[77][23] ), .IN4(n6445), 
        .Q(n2090) );
  AO22X1 U1959 ( .IN1(n6824), .IN2(n6441), .IN3(\FIFO[77][24] ), .IN4(n6446), 
        .Q(n2091) );
  AO22X1 U1960 ( .IN1(n6813), .IN2(n6441), .IN3(\FIFO[77][25] ), .IN4(n6446), 
        .Q(n2092) );
  AO22X1 U1961 ( .IN1(n6802), .IN2(n6441), .IN3(\FIFO[77][26] ), .IN4(n6446), 
        .Q(n2093) );
  AO22X1 U1962 ( .IN1(n6791), .IN2(n6441), .IN3(\FIFO[77][27] ), .IN4(n6446), 
        .Q(n2094) );
  AO22X1 U1963 ( .IN1(n6780), .IN2(n6441), .IN3(\FIFO[77][28] ), .IN4(n6446), 
        .Q(n2095) );
  AO22X1 U1964 ( .IN1(n6769), .IN2(n6442), .IN3(\FIFO[77][29] ), .IN4(n6446), 
        .Q(n2096) );
  AO22X1 U1965 ( .IN1(n6758), .IN2(n6441), .IN3(\FIFO[77][30] ), .IN4(n6446), 
        .Q(n2097) );
  AO22X1 U1966 ( .IN1(n6747), .IN2(n6442), .IN3(\FIFO[77][31] ), .IN4(n6446), 
        .Q(n2098) );
  AO21X1 U1967 ( .IN1(n306), .IN2(n243), .IN3(n7359), .Q(n308) );
  AO22X1 U1968 ( .IN1(n7094), .IN2(n6437), .IN3(\FIFO[76][0] ), .IN4(n6438), 
        .Q(n2099) );
  AO22X1 U1969 ( .IN1(n7077), .IN2(n6436), .IN3(\FIFO[76][1] ), .IN4(n6438), 
        .Q(n2100) );
  AO22X1 U1970 ( .IN1(n7066), .IN2(n6435), .IN3(\FIFO[76][2] ), .IN4(n6438), 
        .Q(n2101) );
  AO22X1 U1971 ( .IN1(n7055), .IN2(n6437), .IN3(\FIFO[76][3] ), .IN4(n6438), 
        .Q(n2102) );
  AO22X1 U1972 ( .IN1(n7044), .IN2(n6436), .IN3(\FIFO[76][4] ), .IN4(n6438), 
        .Q(n2103) );
  AO22X1 U1973 ( .IN1(n7033), .IN2(n6435), .IN3(\FIFO[76][5] ), .IN4(n6438), 
        .Q(n2104) );
  AO22X1 U1974 ( .IN1(n7022), .IN2(n6437), .IN3(\FIFO[76][6] ), .IN4(n6438), 
        .Q(n2105) );
  AO22X1 U1975 ( .IN1(n7011), .IN2(n6437), .IN3(\FIFO[76][7] ), .IN4(n6438), 
        .Q(n2106) );
  AO22X1 U1977 ( .IN1(n6989), .IN2(n6437), .IN3(\FIFO[76][9] ), .IN4(n6438), 
        .Q(n2108) );
  AO22X1 U1978 ( .IN1(n6978), .IN2(n6437), .IN3(\FIFO[76][10] ), .IN4(n6438), 
        .Q(n2109) );
  AO22X1 U1979 ( .IN1(n6967), .IN2(n6437), .IN3(\FIFO[76][11] ), .IN4(n6438), 
        .Q(n2110) );
  AO22X1 U1980 ( .IN1(n6956), .IN2(n6437), .IN3(\FIFO[76][12] ), .IN4(n6439), 
        .Q(n2111) );
  AO22X1 U1981 ( .IN1(n6945), .IN2(n6437), .IN3(\FIFO[76][13] ), .IN4(n6439), 
        .Q(n2112) );
  AO22X1 U1982 ( .IN1(n6934), .IN2(n6436), .IN3(\FIFO[76][14] ), .IN4(n6439), 
        .Q(n2113) );
  AO22X1 U1983 ( .IN1(n6923), .IN2(n6436), .IN3(\FIFO[76][15] ), .IN4(n6439), 
        .Q(n2114) );
  AO22X1 U1984 ( .IN1(n6912), .IN2(n6436), .IN3(\FIFO[76][16] ), .IN4(n6439), 
        .Q(n2115) );
  AO22X1 U1985 ( .IN1(n6901), .IN2(n6436), .IN3(\FIFO[76][17] ), .IN4(n6439), 
        .Q(n2116) );
  AO22X1 U1986 ( .IN1(n6890), .IN2(n6436), .IN3(\FIFO[76][18] ), .IN4(n6439), 
        .Q(n2117) );
  AO22X1 U1987 ( .IN1(n6879), .IN2(n6436), .IN3(\FIFO[76][19] ), .IN4(n6439), 
        .Q(n2118) );
  AO22X1 U1988 ( .IN1(n6868), .IN2(n6436), .IN3(\FIFO[76][20] ), .IN4(n6439), 
        .Q(n2119) );
  AO22X1 U1990 ( .IN1(n6846), .IN2(n6435), .IN3(\FIFO[76][22] ), .IN4(n6439), 
        .Q(n2121) );
  AO22X1 U1991 ( .IN1(n6835), .IN2(n6435), .IN3(\FIFO[76][23] ), .IN4(n6439), 
        .Q(n2122) );
  AO22X1 U1992 ( .IN1(n6824), .IN2(n6435), .IN3(\FIFO[76][24] ), .IN4(n6440), 
        .Q(n2123) );
  AO22X1 U1993 ( .IN1(n6813), .IN2(n6435), .IN3(\FIFO[76][25] ), .IN4(n6440), 
        .Q(n2124) );
  AO22X1 U1994 ( .IN1(n6802), .IN2(n6435), .IN3(\FIFO[76][26] ), .IN4(n6440), 
        .Q(n2125) );
  AO22X1 U1995 ( .IN1(n6791), .IN2(n6435), .IN3(\FIFO[76][27] ), .IN4(n6440), 
        .Q(n2126) );
  AO22X1 U1996 ( .IN1(n6780), .IN2(n6435), .IN3(\FIFO[76][28] ), .IN4(n6440), 
        .Q(n2127) );
  AO22X1 U1997 ( .IN1(n6769), .IN2(n6436), .IN3(\FIFO[76][29] ), .IN4(n6440), 
        .Q(n2128) );
  AO22X1 U1998 ( .IN1(n6758), .IN2(n6435), .IN3(\FIFO[76][30] ), .IN4(n6440), 
        .Q(n2129) );
  AO22X1 U1999 ( .IN1(n6747), .IN2(n6436), .IN3(\FIFO[76][31] ), .IN4(n6440), 
        .Q(n2130) );
  AO21X1 U2000 ( .IN1(n306), .IN2(n245), .IN3(flush), .Q(n309) );
  AO22X1 U2025 ( .IN1(n6824), .IN2(n310), .IN3(\FIFO[75][24] ), .IN4(n6434), 
        .Q(n2155) );
  AO22X1 U2026 ( .IN1(n6813), .IN2(n310), .IN3(\FIFO[75][25] ), .IN4(n6434), 
        .Q(n2156) );
  AO22X1 U2027 ( .IN1(n6802), .IN2(n310), .IN3(\FIFO[75][26] ), .IN4(n6434), 
        .Q(n2157) );
  AO22X1 U2028 ( .IN1(n6791), .IN2(n6431), .IN3(\FIFO[75][27] ), .IN4(n6434), 
        .Q(n2158) );
  AO22X1 U2029 ( .IN1(n6780), .IN2(n6430), .IN3(\FIFO[75][28] ), .IN4(n6434), 
        .Q(n2159) );
  AO22X1 U2030 ( .IN1(n6769), .IN2(n6431), .IN3(\FIFO[75][29] ), .IN4(n6434), 
        .Q(n2160) );
  AO22X1 U2031 ( .IN1(n6758), .IN2(n6430), .IN3(\FIFO[75][30] ), .IN4(n6434), 
        .Q(n2161) );
  AO22X1 U2032 ( .IN1(n6747), .IN2(n6429), .IN3(\FIFO[75][31] ), .IN4(n6434), 
        .Q(n2162) );
  AO21X1 U2033 ( .IN1(n306), .IN2(n247), .IN3(n5973), .Q(n310) );
  AO22X1 U2058 ( .IN1(n6824), .IN2(n311), .IN3(\FIFO[74][24] ), .IN4(n6428), 
        .Q(n2187) );
  AO22X1 U2059 ( .IN1(n6813), .IN2(n311), .IN3(\FIFO[74][25] ), .IN4(n6428), 
        .Q(n2188) );
  AO22X1 U2060 ( .IN1(n6802), .IN2(n311), .IN3(\FIFO[74][26] ), .IN4(n6428), 
        .Q(n2189) );
  AO22X1 U2061 ( .IN1(n6791), .IN2(n6425), .IN3(\FIFO[74][27] ), .IN4(n6428), 
        .Q(n2190) );
  AO22X1 U2062 ( .IN1(n6780), .IN2(n6424), .IN3(\FIFO[74][28] ), .IN4(n6428), 
        .Q(n2191) );
  AO22X1 U2063 ( .IN1(n6769), .IN2(n6425), .IN3(\FIFO[74][29] ), .IN4(n6428), 
        .Q(n2192) );
  AO22X1 U2064 ( .IN1(n6758), .IN2(n6424), .IN3(\FIFO[74][30] ), .IN4(n6428), 
        .Q(n2193) );
  AO22X1 U2065 ( .IN1(n6747), .IN2(n6423), .IN3(\FIFO[74][31] ), .IN4(n6428), 
        .Q(n2194) );
  AO21X1 U2066 ( .IN1(n306), .IN2(n249), .IN3(n7359), .Q(n311) );
  AO22X1 U2067 ( .IN1(n7094), .IN2(n6419), .IN3(\FIFO[73][0] ), .IN4(n6420), 
        .Q(n2195) );
  AO22X1 U2068 ( .IN1(n7077), .IN2(n6419), .IN3(\FIFO[73][1] ), .IN4(n6420), 
        .Q(n2196) );
  AO22X1 U2069 ( .IN1(n7066), .IN2(n6419), .IN3(\FIFO[73][2] ), .IN4(n6420), 
        .Q(n2197) );
  AO22X1 U2070 ( .IN1(n7055), .IN2(n6419), .IN3(\FIFO[73][3] ), .IN4(n6420), 
        .Q(n2198) );
  AO22X1 U2071 ( .IN1(n7044), .IN2(n6419), .IN3(\FIFO[73][4] ), .IN4(n6420), 
        .Q(n2199) );
  AO22X1 U2072 ( .IN1(n7033), .IN2(n6419), .IN3(\FIFO[73][5] ), .IN4(n6420), 
        .Q(n2200) );
  AO22X1 U2073 ( .IN1(n7022), .IN2(n6419), .IN3(\FIFO[73][6] ), .IN4(n6420), 
        .Q(n2201) );
  AO22X1 U2074 ( .IN1(n7011), .IN2(n6418), .IN3(\FIFO[73][7] ), .IN4(n6420), 
        .Q(n2202) );
  AO22X1 U2075 ( .IN1(n7000), .IN2(n6418), .IN3(\FIFO[73][8] ), .IN4(n6420), 
        .Q(n2203) );
  AO22X1 U2076 ( .IN1(n6989), .IN2(n6418), .IN3(\FIFO[73][9] ), .IN4(n6420), 
        .Q(n2204) );
  AO22X1 U2077 ( .IN1(n6978), .IN2(n6418), .IN3(\FIFO[73][10] ), .IN4(n6420), 
        .Q(n2205) );
  AO22X1 U2078 ( .IN1(n6967), .IN2(n6418), .IN3(\FIFO[73][11] ), .IN4(n6420), 
        .Q(n2206) );
  AO22X1 U2079 ( .IN1(n6956), .IN2(n6418), .IN3(\FIFO[73][12] ), .IN4(n6421), 
        .Q(n2207) );
  AO22X1 U2080 ( .IN1(n6945), .IN2(n6418), .IN3(\FIFO[73][13] ), .IN4(n6421), 
        .Q(n2208) );
  AO22X1 U2081 ( .IN1(n6934), .IN2(n6417), .IN3(\FIFO[73][14] ), .IN4(n6421), 
        .Q(n2209) );
  AO22X1 U2082 ( .IN1(n6923), .IN2(n6417), .IN3(\FIFO[73][15] ), .IN4(n6421), 
        .Q(n2210) );
  AO22X1 U2083 ( .IN1(n6912), .IN2(n6417), .IN3(\FIFO[73][16] ), .IN4(n6421), 
        .Q(n2211) );
  AO22X1 U2084 ( .IN1(n6901), .IN2(n6417), .IN3(\FIFO[73][17] ), .IN4(n6421), 
        .Q(n2212) );
  AO22X1 U2085 ( .IN1(n6890), .IN2(n6417), .IN3(\FIFO[73][18] ), .IN4(n6421), 
        .Q(n2213) );
  AO22X1 U2086 ( .IN1(n6879), .IN2(n6417), .IN3(\FIFO[73][19] ), .IN4(n6421), 
        .Q(n2214) );
  AO22X1 U2087 ( .IN1(n6868), .IN2(n6417), .IN3(\FIFO[73][20] ), .IN4(n6421), 
        .Q(n2215) );
  AO22X1 U2088 ( .IN1(n6857), .IN2(n6419), .IN3(\FIFO[73][21] ), .IN4(n6421), 
        .Q(n2216) );
  AO22X1 U2089 ( .IN1(n6846), .IN2(n6418), .IN3(\FIFO[73][22] ), .IN4(n6421), 
        .Q(n2217) );
  AO22X1 U2090 ( .IN1(n6835), .IN2(n6417), .IN3(\FIFO[73][23] ), .IN4(n6421), 
        .Q(n2218) );
  AO22X1 U2091 ( .IN1(n6824), .IN2(n312), .IN3(\FIFO[73][24] ), .IN4(n6422), 
        .Q(n2219) );
  AO22X1 U2092 ( .IN1(n6813), .IN2(n312), .IN3(\FIFO[73][25] ), .IN4(n6422), 
        .Q(n2220) );
  AO22X1 U2093 ( .IN1(n6802), .IN2(n312), .IN3(\FIFO[73][26] ), .IN4(n6422), 
        .Q(n2221) );
  AO22X1 U2094 ( .IN1(n6791), .IN2(n6419), .IN3(\FIFO[73][27] ), .IN4(n6422), 
        .Q(n2222) );
  AO22X1 U2095 ( .IN1(n6780), .IN2(n6419), .IN3(\FIFO[73][28] ), .IN4(n6422), 
        .Q(n2223) );
  AO22X1 U2096 ( .IN1(n6769), .IN2(n6418), .IN3(\FIFO[73][29] ), .IN4(n6422), 
        .Q(n2224) );
  AO22X1 U2097 ( .IN1(n6758), .IN2(n6417), .IN3(\FIFO[73][30] ), .IN4(n6422), 
        .Q(n2225) );
  AO22X1 U2098 ( .IN1(n6747), .IN2(n6418), .IN3(\FIFO[73][31] ), .IN4(n6422), 
        .Q(n2226) );
  AO21X1 U2099 ( .IN1(n306), .IN2(n251), .IN3(flush), .Q(n312) );
  AO22X1 U2100 ( .IN1(n7094), .IN2(n6413), .IN3(\FIFO[72][0] ), .IN4(n6414), 
        .Q(n2227) );
  AO22X1 U2101 ( .IN1(n7077), .IN2(n6413), .IN3(\FIFO[72][1] ), .IN4(n6414), 
        .Q(n2228) );
  AO22X1 U2102 ( .IN1(n7066), .IN2(n6413), .IN3(\FIFO[72][2] ), .IN4(n6414), 
        .Q(n2229) );
  AO22X1 U2103 ( .IN1(n7055), .IN2(n6413), .IN3(\FIFO[72][3] ), .IN4(n6414), 
        .Q(n2230) );
  AO22X1 U2104 ( .IN1(n7044), .IN2(n6413), .IN3(\FIFO[72][4] ), .IN4(n6414), 
        .Q(n2231) );
  AO22X1 U2105 ( .IN1(n7033), .IN2(n6413), .IN3(\FIFO[72][5] ), .IN4(n6414), 
        .Q(n2232) );
  AO22X1 U2106 ( .IN1(n7022), .IN2(n6413), .IN3(\FIFO[72][6] ), .IN4(n6414), 
        .Q(n2233) );
  AO22X1 U2107 ( .IN1(n7011), .IN2(n6412), .IN3(\FIFO[72][7] ), .IN4(n6414), 
        .Q(n2234) );
  AO22X1 U2108 ( .IN1(n7000), .IN2(n6412), .IN3(\FIFO[72][8] ), .IN4(n6414), 
        .Q(n2235) );
  AO22X1 U2110 ( .IN1(n6978), .IN2(n6412), .IN3(\FIFO[72][10] ), .IN4(n6414), 
        .Q(n2237) );
  AO22X1 U2111 ( .IN1(n6967), .IN2(n6412), .IN3(\FIFO[72][11] ), .IN4(n6414), 
        .Q(n2238) );
  AO22X1 U2112 ( .IN1(n6956), .IN2(n6412), .IN3(\FIFO[72][12] ), .IN4(n6415), 
        .Q(n2239) );
  AO22X1 U2113 ( .IN1(n6945), .IN2(n6412), .IN3(\FIFO[72][13] ), .IN4(n6415), 
        .Q(n2240) );
  AO22X1 U2114 ( .IN1(n6934), .IN2(n6413), .IN3(\FIFO[72][14] ), .IN4(n6415), 
        .Q(n2241) );
  AO22X1 U2115 ( .IN1(n6923), .IN2(n6412), .IN3(\FIFO[72][15] ), .IN4(n6415), 
        .Q(n2242) );
  AO22X1 U2116 ( .IN1(n6912), .IN2(n6411), .IN3(\FIFO[72][16] ), .IN4(n6415), 
        .Q(n2243) );
  AO22X1 U2117 ( .IN1(n6901), .IN2(n6413), .IN3(\FIFO[72][17] ), .IN4(n6415), 
        .Q(n2244) );
  AO22X1 U2118 ( .IN1(n6890), .IN2(n6412), .IN3(\FIFO[72][18] ), .IN4(n6415), 
        .Q(n2245) );
  AO22X1 U2119 ( .IN1(n6879), .IN2(n6411), .IN3(\FIFO[72][19] ), .IN4(n6415), 
        .Q(n2246) );
  AO22X1 U2120 ( .IN1(n6868), .IN2(n6413), .IN3(\FIFO[72][20] ), .IN4(n6415), 
        .Q(n2247) );
  AO22X1 U2121 ( .IN1(n6857), .IN2(n6411), .IN3(\FIFO[72][21] ), .IN4(n6415), 
        .Q(n2248) );
  AO22X1 U2123 ( .IN1(n6835), .IN2(n6411), .IN3(\FIFO[72][23] ), .IN4(n6415), 
        .Q(n2250) );
  AO22X1 U2124 ( .IN1(n6824), .IN2(n6411), .IN3(\FIFO[72][24] ), .IN4(n6416), 
        .Q(n2251) );
  AO22X1 U2125 ( .IN1(n6813), .IN2(n6411), .IN3(\FIFO[72][25] ), .IN4(n6416), 
        .Q(n2252) );
  AO22X1 U2126 ( .IN1(n6802), .IN2(n6411), .IN3(\FIFO[72][26] ), .IN4(n6416), 
        .Q(n2253) );
  AO22X1 U2127 ( .IN1(n6791), .IN2(n6411), .IN3(\FIFO[72][27] ), .IN4(n6416), 
        .Q(n2254) );
  AO22X1 U2128 ( .IN1(n6780), .IN2(n6411), .IN3(\FIFO[72][28] ), .IN4(n6416), 
        .Q(n2255) );
  AO22X1 U2129 ( .IN1(n6769), .IN2(n6412), .IN3(\FIFO[72][29] ), .IN4(n6416), 
        .Q(n2256) );
  AO22X1 U2130 ( .IN1(n6758), .IN2(n6411), .IN3(\FIFO[72][30] ), .IN4(n6416), 
        .Q(n2257) );
  AO22X1 U2131 ( .IN1(n6747), .IN2(n6412), .IN3(\FIFO[72][31] ), .IN4(n6416), 
        .Q(n2258) );
  AO21X1 U2132 ( .IN1(n306), .IN2(n253), .IN3(n5973), .Q(n313) );
  AO22X1 U2157 ( .IN1(n6823), .IN2(n6405), .IN3(\FIFO[71][24] ), .IN4(n6410), 
        .Q(n2283) );
  AO22X1 U2158 ( .IN1(n6812), .IN2(n6405), .IN3(\FIFO[71][25] ), .IN4(n6410), 
        .Q(n2284) );
  AO22X1 U2159 ( .IN1(n6801), .IN2(n6405), .IN3(\FIFO[71][26] ), .IN4(n6410), 
        .Q(n2285) );
  AO22X1 U2160 ( .IN1(n6790), .IN2(n6405), .IN3(\FIFO[71][27] ), .IN4(n6410), 
        .Q(n2286) );
  AO22X1 U2161 ( .IN1(n6779), .IN2(n6405), .IN3(\FIFO[71][28] ), .IN4(n6410), 
        .Q(n2287) );
  AO22X1 U2162 ( .IN1(n6768), .IN2(n6406), .IN3(\FIFO[71][29] ), .IN4(n6410), 
        .Q(n2288) );
  AO22X1 U2163 ( .IN1(n6757), .IN2(n6405), .IN3(\FIFO[71][30] ), .IN4(n6410), 
        .Q(n2289) );
  AO22X1 U2164 ( .IN1(n6746), .IN2(n6406), .IN3(\FIFO[71][31] ), .IN4(n6410), 
        .Q(n2290) );
  AO21X1 U2165 ( .IN1(n306), .IN2(n255), .IN3(n7359), .Q(n314) );
  AO22X1 U2190 ( .IN1(n6823), .IN2(n315), .IN3(\FIFO[70][24] ), .IN4(n6404), 
        .Q(n2315) );
  AO22X1 U2191 ( .IN1(n6812), .IN2(n315), .IN3(\FIFO[70][25] ), .IN4(n6404), 
        .Q(n2316) );
  AO22X1 U2192 ( .IN1(n6801), .IN2(n315), .IN3(\FIFO[70][26] ), .IN4(n6404), 
        .Q(n2317) );
  AO22X1 U2193 ( .IN1(n6790), .IN2(n6401), .IN3(\FIFO[70][27] ), .IN4(n6404), 
        .Q(n2318) );
  AO22X1 U2194 ( .IN1(n6779), .IN2(n6400), .IN3(\FIFO[70][28] ), .IN4(n6404), 
        .Q(n2319) );
  AO22X1 U2195 ( .IN1(n6768), .IN2(n6401), .IN3(\FIFO[70][29] ), .IN4(n6404), 
        .Q(n2320) );
  AO22X1 U2196 ( .IN1(n6757), .IN2(n6400), .IN3(\FIFO[70][30] ), .IN4(n6404), 
        .Q(n2321) );
  AO22X1 U2197 ( .IN1(n6746), .IN2(n6399), .IN3(\FIFO[70][31] ), .IN4(n6404), 
        .Q(n2322) );
  AO21X1 U2198 ( .IN1(n306), .IN2(n257), .IN3(flush), .Q(n315) );
  AO22X1 U2199 ( .IN1(n7093), .IN2(n6395), .IN3(\FIFO[69][0] ), .IN4(n6396), 
        .Q(n2323) );
  AO22X1 U2200 ( .IN1(n7076), .IN2(n6395), .IN3(\FIFO[69][1] ), .IN4(n6396), 
        .Q(n2324) );
  AO22X1 U2201 ( .IN1(n7065), .IN2(n6395), .IN3(\FIFO[69][2] ), .IN4(n6396), 
        .Q(n2325) );
  AO22X1 U2202 ( .IN1(n7054), .IN2(n6395), .IN3(\FIFO[69][3] ), .IN4(n6396), 
        .Q(n2326) );
  AO22X1 U2203 ( .IN1(n7043), .IN2(n6395), .IN3(\FIFO[69][4] ), .IN4(n6396), 
        .Q(n2327) );
  AO22X1 U2204 ( .IN1(n7032), .IN2(n6395), .IN3(\FIFO[69][5] ), .IN4(n6396), 
        .Q(n2328) );
  AO22X1 U2205 ( .IN1(n7021), .IN2(n6395), .IN3(\FIFO[69][6] ), .IN4(n6396), 
        .Q(n2329) );
  AO22X1 U2206 ( .IN1(n7010), .IN2(n6394), .IN3(\FIFO[69][7] ), .IN4(n6396), 
        .Q(n2330) );
  AO22X1 U2207 ( .IN1(n6999), .IN2(n6394), .IN3(\FIFO[69][8] ), .IN4(n6396), 
        .Q(n2331) );
  AO22X1 U2208 ( .IN1(n6988), .IN2(n6394), .IN3(\FIFO[69][9] ), .IN4(n6396), 
        .Q(n2332) );
  AO22X1 U2209 ( .IN1(n6977), .IN2(n6394), .IN3(\FIFO[69][10] ), .IN4(n6396), 
        .Q(n2333) );
  AO22X1 U2210 ( .IN1(n6966), .IN2(n6394), .IN3(\FIFO[69][11] ), .IN4(n6396), 
        .Q(n2334) );
  AO22X1 U2211 ( .IN1(n6955), .IN2(n6394), .IN3(\FIFO[69][12] ), .IN4(n6397), 
        .Q(n2335) );
  AO22X1 U2212 ( .IN1(n6944), .IN2(n6394), .IN3(\FIFO[69][13] ), .IN4(n6397), 
        .Q(n2336) );
  AO22X1 U2213 ( .IN1(n6933), .IN2(n6393), .IN3(\FIFO[69][14] ), .IN4(n6397), 
        .Q(n2337) );
  AO22X1 U2214 ( .IN1(n6922), .IN2(n6393), .IN3(\FIFO[69][15] ), .IN4(n6397), 
        .Q(n2338) );
  AO22X1 U2215 ( .IN1(n6911), .IN2(n6393), .IN3(\FIFO[69][16] ), .IN4(n6397), 
        .Q(n2339) );
  AO22X1 U2216 ( .IN1(n6900), .IN2(n6393), .IN3(\FIFO[69][17] ), .IN4(n6397), 
        .Q(n2340) );
  AO22X1 U2217 ( .IN1(n6889), .IN2(n6393), .IN3(\FIFO[69][18] ), .IN4(n6397), 
        .Q(n2341) );
  AO22X1 U2218 ( .IN1(n6878), .IN2(n6393), .IN3(\FIFO[69][19] ), .IN4(n6397), 
        .Q(n2342) );
  AO22X1 U2219 ( .IN1(n6867), .IN2(n6393), .IN3(\FIFO[69][20] ), .IN4(n6397), 
        .Q(n2343) );
  AO22X1 U2220 ( .IN1(n6856), .IN2(n6395), .IN3(\FIFO[69][21] ), .IN4(n6397), 
        .Q(n2344) );
  AO22X1 U2221 ( .IN1(n6845), .IN2(n6394), .IN3(\FIFO[69][22] ), .IN4(n6397), 
        .Q(n2345) );
  AO22X1 U2222 ( .IN1(n6834), .IN2(n6393), .IN3(\FIFO[69][23] ), .IN4(n6397), 
        .Q(n2346) );
  AO22X1 U2223 ( .IN1(n6823), .IN2(n316), .IN3(\FIFO[69][24] ), .IN4(n6398), 
        .Q(n2347) );
  AO22X1 U2224 ( .IN1(n6812), .IN2(n316), .IN3(\FIFO[69][25] ), .IN4(n6398), 
        .Q(n2348) );
  AO22X1 U2225 ( .IN1(n6801), .IN2(n316), .IN3(\FIFO[69][26] ), .IN4(n6398), 
        .Q(n2349) );
  AO22X1 U2226 ( .IN1(n6790), .IN2(n6395), .IN3(\FIFO[69][27] ), .IN4(n6398), 
        .Q(n2350) );
  AO22X1 U2227 ( .IN1(n6779), .IN2(n6394), .IN3(\FIFO[69][28] ), .IN4(n6398), 
        .Q(n2351) );
  AO22X1 U2228 ( .IN1(n6768), .IN2(n6395), .IN3(\FIFO[69][29] ), .IN4(n6398), 
        .Q(n2352) );
  AO22X1 U2229 ( .IN1(n6757), .IN2(n6394), .IN3(\FIFO[69][30] ), .IN4(n6398), 
        .Q(n2353) );
  AO22X1 U2230 ( .IN1(n6746), .IN2(n6393), .IN3(\FIFO[69][31] ), .IN4(n6398), 
        .Q(n2354) );
  AO21X1 U2231 ( .IN1(n306), .IN2(n259), .IN3(n5973), .Q(n316) );
  AO22X1 U2232 ( .IN1(n7093), .IN2(n6389), .IN3(\FIFO[68][0] ), .IN4(n6390), 
        .Q(n2355) );
  AO22X1 U2233 ( .IN1(n7076), .IN2(n6389), .IN3(\FIFO[68][1] ), .IN4(n6390), 
        .Q(n2356) );
  AO22X1 U2234 ( .IN1(n7065), .IN2(n6389), .IN3(\FIFO[68][2] ), .IN4(n6390), 
        .Q(n2357) );
  AO22X1 U2235 ( .IN1(n7054), .IN2(n6389), .IN3(\FIFO[68][3] ), .IN4(n6390), 
        .Q(n2358) );
  AO22X1 U2236 ( .IN1(n7043), .IN2(n6389), .IN3(\FIFO[68][4] ), .IN4(n6390), 
        .Q(n2359) );
  AO22X1 U2237 ( .IN1(n7032), .IN2(n6389), .IN3(\FIFO[68][5] ), .IN4(n6390), 
        .Q(n2360) );
  AO22X1 U2238 ( .IN1(n7021), .IN2(n6389), .IN3(\FIFO[68][6] ), .IN4(n6390), 
        .Q(n2361) );
  AO22X1 U2239 ( .IN1(n7010), .IN2(n6388), .IN3(\FIFO[68][7] ), .IN4(n6390), 
        .Q(n2362) );
  AO22X1 U2240 ( .IN1(n6999), .IN2(n6388), .IN3(\FIFO[68][8] ), .IN4(n6390), 
        .Q(n2363) );
  AO22X1 U2241 ( .IN1(n6988), .IN2(n6388), .IN3(\FIFO[68][9] ), .IN4(n6390), 
        .Q(n2364) );
  AO22X1 U2242 ( .IN1(n6977), .IN2(n6388), .IN3(\FIFO[68][10] ), .IN4(n6390), 
        .Q(n2365) );
  AO22X1 U2243 ( .IN1(n6966), .IN2(n6388), .IN3(\FIFO[68][11] ), .IN4(n6390), 
        .Q(n2366) );
  AO22X1 U2244 ( .IN1(n6955), .IN2(n6388), .IN3(\FIFO[68][12] ), .IN4(n6391), 
        .Q(n2367) );
  AO22X1 U2245 ( .IN1(n6944), .IN2(n6388), .IN3(\FIFO[68][13] ), .IN4(n6391), 
        .Q(n2368) );
  AO22X1 U2246 ( .IN1(n6933), .IN2(n6387), .IN3(\FIFO[68][14] ), .IN4(n6391), 
        .Q(n2369) );
  AO22X1 U2247 ( .IN1(n6922), .IN2(n6387), .IN3(\FIFO[68][15] ), .IN4(n6391), 
        .Q(n2370) );
  AO22X1 U2248 ( .IN1(n6911), .IN2(n6387), .IN3(\FIFO[68][16] ), .IN4(n6391), 
        .Q(n2371) );
  AO22X1 U2249 ( .IN1(n6900), .IN2(n6387), .IN3(\FIFO[68][17] ), .IN4(n6391), 
        .Q(n2372) );
  AO22X1 U2250 ( .IN1(n6889), .IN2(n6387), .IN3(\FIFO[68][18] ), .IN4(n6391), 
        .Q(n2373) );
  AO22X1 U2251 ( .IN1(n6878), .IN2(n6387), .IN3(\FIFO[68][19] ), .IN4(n6391), 
        .Q(n2374) );
  AO22X1 U2252 ( .IN1(n6867), .IN2(n6387), .IN3(\FIFO[68][20] ), .IN4(n6391), 
        .Q(n2375) );
  AO22X1 U2253 ( .IN1(n6856), .IN2(n6389), .IN3(\FIFO[68][21] ), .IN4(n6391), 
        .Q(n2376) );
  AO22X1 U2254 ( .IN1(n6845), .IN2(n6388), .IN3(\FIFO[68][22] ), .IN4(n6391), 
        .Q(n2377) );
  AO22X1 U2255 ( .IN1(n6834), .IN2(n6387), .IN3(\FIFO[68][23] ), .IN4(n6391), 
        .Q(n2378) );
  AO22X1 U2256 ( .IN1(n6823), .IN2(n317), .IN3(\FIFO[68][24] ), .IN4(n6392), 
        .Q(n2379) );
  AO22X1 U2257 ( .IN1(n6812), .IN2(n317), .IN3(\FIFO[68][25] ), .IN4(n6392), 
        .Q(n2380) );
  AO22X1 U2258 ( .IN1(n6801), .IN2(n317), .IN3(\FIFO[68][26] ), .IN4(n6392), 
        .Q(n2381) );
  AO22X1 U2259 ( .IN1(n6790), .IN2(n6389), .IN3(\FIFO[68][27] ), .IN4(n6392), 
        .Q(n2382) );
  AO22X1 U2260 ( .IN1(n6779), .IN2(n6389), .IN3(\FIFO[68][28] ), .IN4(n6392), 
        .Q(n2383) );
  AO22X1 U2261 ( .IN1(n6768), .IN2(n6388), .IN3(\FIFO[68][29] ), .IN4(n6392), 
        .Q(n2384) );
  AO22X1 U2262 ( .IN1(n6757), .IN2(n6387), .IN3(\FIFO[68][30] ), .IN4(n6392), 
        .Q(n2385) );
  AO22X1 U2263 ( .IN1(n6746), .IN2(n6388), .IN3(\FIFO[68][31] ), .IN4(n6392), 
        .Q(n2386) );
  AO21X1 U2264 ( .IN1(n306), .IN2(n261), .IN3(n7359), .Q(n317) );
  AO22X1 U2289 ( .IN1(n6823), .IN2(n6381), .IN3(\FIFO[67][24] ), .IN4(n6386), 
        .Q(n2411) );
  AO22X1 U2290 ( .IN1(n6812), .IN2(n6381), .IN3(\FIFO[67][25] ), .IN4(n6386), 
        .Q(n2412) );
  AO22X1 U2291 ( .IN1(n6801), .IN2(n6381), .IN3(\FIFO[67][26] ), .IN4(n6386), 
        .Q(n2413) );
  AO22X1 U2292 ( .IN1(n6790), .IN2(n6381), .IN3(\FIFO[67][27] ), .IN4(n6386), 
        .Q(n2414) );
  AO22X1 U2293 ( .IN1(n6779), .IN2(n6381), .IN3(\FIFO[67][28] ), .IN4(n6386), 
        .Q(n2415) );
  AO22X1 U2294 ( .IN1(n6768), .IN2(n6382), .IN3(\FIFO[67][29] ), .IN4(n6386), 
        .Q(n2416) );
  AO22X1 U2295 ( .IN1(n6757), .IN2(n6381), .IN3(\FIFO[67][30] ), .IN4(n6386), 
        .Q(n2417) );
  AO22X1 U2296 ( .IN1(n6746), .IN2(n6382), .IN3(\FIFO[67][31] ), .IN4(n6386), 
        .Q(n2418) );
  AO21X1 U2297 ( .IN1(n306), .IN2(n263), .IN3(flush), .Q(n318) );
  AO22X1 U2322 ( .IN1(n6823), .IN2(n6375), .IN3(\FIFO[66][24] ), .IN4(n6380), 
        .Q(n2443) );
  AO22X1 U2323 ( .IN1(n6812), .IN2(n6375), .IN3(\FIFO[66][25] ), .IN4(n6380), 
        .Q(n2444) );
  AO22X1 U2324 ( .IN1(n6801), .IN2(n6375), .IN3(\FIFO[66][26] ), .IN4(n6380), 
        .Q(n2445) );
  AO22X1 U2325 ( .IN1(n6790), .IN2(n6375), .IN3(\FIFO[66][27] ), .IN4(n6380), 
        .Q(n2446) );
  AO22X1 U2326 ( .IN1(n6779), .IN2(n6375), .IN3(\FIFO[66][28] ), .IN4(n6380), 
        .Q(n2447) );
  AO22X1 U2327 ( .IN1(n6768), .IN2(n6376), .IN3(\FIFO[66][29] ), .IN4(n6380), 
        .Q(n2448) );
  AO22X1 U2328 ( .IN1(n6757), .IN2(n6375), .IN3(\FIFO[66][30] ), .IN4(n6380), 
        .Q(n2449) );
  AO22X1 U2329 ( .IN1(n6746), .IN2(n6376), .IN3(\FIFO[66][31] ), .IN4(n6380), 
        .Q(n2450) );
  AO21X1 U2330 ( .IN1(n306), .IN2(n265), .IN3(n5973), .Q(n319) );
  AO22X1 U2331 ( .IN1(n7093), .IN2(n6371), .IN3(\FIFO[65][0] ), .IN4(n6372), 
        .Q(n2451) );
  AO22X1 U2332 ( .IN1(n7076), .IN2(n6371), .IN3(\FIFO[65][1] ), .IN4(n6372), 
        .Q(n2452) );
  AO22X1 U2333 ( .IN1(n7065), .IN2(n6371), .IN3(\FIFO[65][2] ), .IN4(n6372), 
        .Q(n2453) );
  AO22X1 U2334 ( .IN1(n7054), .IN2(n6371), .IN3(\FIFO[65][3] ), .IN4(n6372), 
        .Q(n2454) );
  AO22X1 U2335 ( .IN1(n7043), .IN2(n6371), .IN3(\FIFO[65][4] ), .IN4(n6372), 
        .Q(n2455) );
  AO22X1 U2336 ( .IN1(n7032), .IN2(n6371), .IN3(\FIFO[65][5] ), .IN4(n6372), 
        .Q(n2456) );
  AO22X1 U2337 ( .IN1(n7021), .IN2(n6371), .IN3(\FIFO[65][6] ), .IN4(n6372), 
        .Q(n2457) );
  AO22X1 U2338 ( .IN1(n7010), .IN2(n6370), .IN3(\FIFO[65][7] ), .IN4(n6372), 
        .Q(n2458) );
  AO22X1 U2339 ( .IN1(n6999), .IN2(n6370), .IN3(\FIFO[65][8] ), .IN4(n6372), 
        .Q(n2459) );
  AO22X1 U2340 ( .IN1(n6988), .IN2(n6370), .IN3(\FIFO[65][9] ), .IN4(n6372), 
        .Q(n2460) );
  AO22X1 U2341 ( .IN1(n6977), .IN2(n6370), .IN3(\FIFO[65][10] ), .IN4(n6372), 
        .Q(n2461) );
  AO22X1 U2342 ( .IN1(n6966), .IN2(n6370), .IN3(\FIFO[65][11] ), .IN4(n6372), 
        .Q(n2462) );
  AO22X1 U2343 ( .IN1(n6955), .IN2(n6370), .IN3(\FIFO[65][12] ), .IN4(n6373), 
        .Q(n2463) );
  AO22X1 U2344 ( .IN1(n6944), .IN2(n6370), .IN3(\FIFO[65][13] ), .IN4(n6373), 
        .Q(n2464) );
  AO22X1 U2345 ( .IN1(n6933), .IN2(n6369), .IN3(\FIFO[65][14] ), .IN4(n6373), 
        .Q(n2465) );
  AO22X1 U2346 ( .IN1(n6922), .IN2(n6369), .IN3(\FIFO[65][15] ), .IN4(n6373), 
        .Q(n2466) );
  AO22X1 U2347 ( .IN1(n6911), .IN2(n6369), .IN3(\FIFO[65][16] ), .IN4(n6373), 
        .Q(n2467) );
  AO22X1 U2348 ( .IN1(n6900), .IN2(n6369), .IN3(\FIFO[65][17] ), .IN4(n6373), 
        .Q(n2468) );
  AO22X1 U2349 ( .IN1(n6889), .IN2(n6369), .IN3(\FIFO[65][18] ), .IN4(n6373), 
        .Q(n2469) );
  AO22X1 U2350 ( .IN1(n6878), .IN2(n6369), .IN3(\FIFO[65][19] ), .IN4(n6373), 
        .Q(n2470) );
  AO22X1 U2351 ( .IN1(n6867), .IN2(n6369), .IN3(\FIFO[65][20] ), .IN4(n6373), 
        .Q(n2471) );
  AO22X1 U2352 ( .IN1(n6856), .IN2(n6371), .IN3(\FIFO[65][21] ), .IN4(n6373), 
        .Q(n2472) );
  AO22X1 U2353 ( .IN1(n6845), .IN2(n6370), .IN3(\FIFO[65][22] ), .IN4(n6373), 
        .Q(n2473) );
  AO22X1 U2354 ( .IN1(n6834), .IN2(n6369), .IN3(\FIFO[65][23] ), .IN4(n6373), 
        .Q(n2474) );
  AO22X1 U2355 ( .IN1(n6823), .IN2(n320), .IN3(\FIFO[65][24] ), .IN4(n6374), 
        .Q(n2475) );
  AO22X1 U2356 ( .IN1(n6812), .IN2(n320), .IN3(\FIFO[65][25] ), .IN4(n6374), 
        .Q(n2476) );
  AO22X1 U2357 ( .IN1(n6801), .IN2(n320), .IN3(\FIFO[65][26] ), .IN4(n6374), 
        .Q(n2477) );
  AO22X1 U2358 ( .IN1(n6790), .IN2(n6371), .IN3(\FIFO[65][27] ), .IN4(n6374), 
        .Q(n2478) );
  AO22X1 U2359 ( .IN1(n6779), .IN2(n6370), .IN3(\FIFO[65][28] ), .IN4(n6374), 
        .Q(n2479) );
  AO22X1 U2360 ( .IN1(n6768), .IN2(n6371), .IN3(\FIFO[65][29] ), .IN4(n6374), 
        .Q(n2480) );
  AO22X1 U2361 ( .IN1(n6757), .IN2(n6370), .IN3(\FIFO[65][30] ), .IN4(n6374), 
        .Q(n2481) );
  AO22X1 U2362 ( .IN1(n6746), .IN2(n6369), .IN3(\FIFO[65][31] ), .IN4(n6374), 
        .Q(n2482) );
  AO21X1 U2363 ( .IN1(n306), .IN2(n267), .IN3(n7359), .Q(n320) );
  AO22X1 U2364 ( .IN1(n7093), .IN2(n6365), .IN3(\FIFO[64][0] ), .IN4(n6366), 
        .Q(n2483) );
  AO22X1 U2365 ( .IN1(n7076), .IN2(n6365), .IN3(\FIFO[64][1] ), .IN4(n6366), 
        .Q(n2484) );
  AO22X1 U2366 ( .IN1(n7065), .IN2(n6365), .IN3(\FIFO[64][2] ), .IN4(n6366), 
        .Q(n2485) );
  AO22X1 U2367 ( .IN1(n7054), .IN2(n6365), .IN3(\FIFO[64][3] ), .IN4(n6366), 
        .Q(n2486) );
  AO22X1 U2368 ( .IN1(n7043), .IN2(n6365), .IN3(\FIFO[64][4] ), .IN4(n6366), 
        .Q(n2487) );
  AO22X1 U2369 ( .IN1(n7032), .IN2(n6365), .IN3(\FIFO[64][5] ), .IN4(n6366), 
        .Q(n2488) );
  AO22X1 U2370 ( .IN1(n7021), .IN2(n6365), .IN3(\FIFO[64][6] ), .IN4(n6366), 
        .Q(n2489) );
  AO22X1 U2371 ( .IN1(n7010), .IN2(n6364), .IN3(\FIFO[64][7] ), .IN4(n6366), 
        .Q(n2490) );
  AO22X1 U2372 ( .IN1(n6999), .IN2(n6364), .IN3(\FIFO[64][8] ), .IN4(n6366), 
        .Q(n2491) );
  AO22X1 U2373 ( .IN1(n6988), .IN2(n6364), .IN3(\FIFO[64][9] ), .IN4(n6366), 
        .Q(n2492) );
  AO22X1 U2374 ( .IN1(n6977), .IN2(n6364), .IN3(\FIFO[64][10] ), .IN4(n6366), 
        .Q(n2493) );
  AO22X1 U2375 ( .IN1(n6966), .IN2(n6364), .IN3(\FIFO[64][11] ), .IN4(n6366), 
        .Q(n2494) );
  AO22X1 U2376 ( .IN1(n6955), .IN2(n6364), .IN3(\FIFO[64][12] ), .IN4(n6367), 
        .Q(n2495) );
  AO22X1 U2377 ( .IN1(n6944), .IN2(n6364), .IN3(\FIFO[64][13] ), .IN4(n6367), 
        .Q(n2496) );
  AO22X1 U2378 ( .IN1(n6933), .IN2(n6363), .IN3(\FIFO[64][14] ), .IN4(n6367), 
        .Q(n2497) );
  AO22X1 U2379 ( .IN1(n6922), .IN2(n6363), .IN3(\FIFO[64][15] ), .IN4(n6367), 
        .Q(n2498) );
  AO22X1 U2380 ( .IN1(n6911), .IN2(n6363), .IN3(\FIFO[64][16] ), .IN4(n6367), 
        .Q(n2499) );
  AO22X1 U2381 ( .IN1(n6900), .IN2(n6363), .IN3(\FIFO[64][17] ), .IN4(n6367), 
        .Q(n2500) );
  AO22X1 U2382 ( .IN1(n6889), .IN2(n6363), .IN3(\FIFO[64][18] ), .IN4(n6367), 
        .Q(n2501) );
  AO22X1 U2383 ( .IN1(n6878), .IN2(n6363), .IN3(\FIFO[64][19] ), .IN4(n6367), 
        .Q(n2502) );
  AO22X1 U2384 ( .IN1(n6867), .IN2(n6363), .IN3(\FIFO[64][20] ), .IN4(n6367), 
        .Q(n2503) );
  AO22X1 U2385 ( .IN1(n6856), .IN2(n6365), .IN3(\FIFO[64][21] ), .IN4(n6367), 
        .Q(n2504) );
  AO22X1 U2386 ( .IN1(n6845), .IN2(n6364), .IN3(\FIFO[64][22] ), .IN4(n6367), 
        .Q(n2505) );
  AO22X1 U2387 ( .IN1(n6834), .IN2(n6363), .IN3(\FIFO[64][23] ), .IN4(n6367), 
        .Q(n2506) );
  AO22X1 U2388 ( .IN1(n6823), .IN2(n321), .IN3(\FIFO[64][24] ), .IN4(n6368), 
        .Q(n2507) );
  AO22X1 U2389 ( .IN1(n6812), .IN2(n321), .IN3(\FIFO[64][25] ), .IN4(n6368), 
        .Q(n2508) );
  AO22X1 U2390 ( .IN1(n6801), .IN2(n321), .IN3(\FIFO[64][26] ), .IN4(n6368), 
        .Q(n2509) );
  AO22X1 U2391 ( .IN1(n6790), .IN2(n6365), .IN3(\FIFO[64][27] ), .IN4(n6368), 
        .Q(n2510) );
  AO22X1 U2392 ( .IN1(n6779), .IN2(n6364), .IN3(\FIFO[64][28] ), .IN4(n6368), 
        .Q(n2511) );
  AO22X1 U2393 ( .IN1(n6768), .IN2(n6365), .IN3(\FIFO[64][29] ), .IN4(n6368), 
        .Q(n2512) );
  AO22X1 U2394 ( .IN1(n6757), .IN2(n6364), .IN3(\FIFO[64][30] ), .IN4(n6368), 
        .Q(n2513) );
  AO22X1 U2395 ( .IN1(n6746), .IN2(n6363), .IN3(\FIFO[64][31] ), .IN4(n6368), 
        .Q(n2514) );
  AO21X1 U2396 ( .IN1(n306), .IN2(n269), .IN3(n5973), .Q(n321) );
  AO22X1 U2422 ( .IN1(n6823), .IN2(n6357), .IN3(\FIFO[63][24] ), .IN4(n6362), 
        .Q(n2539) );
  AO22X1 U2423 ( .IN1(n6812), .IN2(n6357), .IN3(\FIFO[63][25] ), .IN4(n6362), 
        .Q(n2540) );
  AO22X1 U2424 ( .IN1(n6801), .IN2(n6357), .IN3(\FIFO[63][26] ), .IN4(n6362), 
        .Q(n2541) );
  AO22X1 U2425 ( .IN1(n6790), .IN2(n6357), .IN3(\FIFO[63][27] ), .IN4(n6362), 
        .Q(n2542) );
  AO22X1 U2426 ( .IN1(n6779), .IN2(n6357), .IN3(\FIFO[63][28] ), .IN4(n6362), 
        .Q(n2543) );
  AO22X1 U2427 ( .IN1(n6768), .IN2(n6358), .IN3(\FIFO[63][29] ), .IN4(n6362), 
        .Q(n2544) );
  AO22X1 U2428 ( .IN1(n6757), .IN2(n6357), .IN3(\FIFO[63][30] ), .IN4(n6362), 
        .Q(n2545) );
  AO22X1 U2429 ( .IN1(n6746), .IN2(n6358), .IN3(\FIFO[63][31] ), .IN4(n6362), 
        .Q(n2546) );
  AO21X1 U2430 ( .IN1(n323), .IN2(n238), .IN3(n7359), .Q(n322) );
  AO22X1 U2455 ( .IN1(n6823), .IN2(n6351), .IN3(\FIFO[62][24] ), .IN4(n6356), 
        .Q(n2571) );
  AO22X1 U2456 ( .IN1(n6812), .IN2(n6351), .IN3(\FIFO[62][25] ), .IN4(n6356), 
        .Q(n2572) );
  AO22X1 U2457 ( .IN1(n6801), .IN2(n6351), .IN3(\FIFO[62][26] ), .IN4(n6356), 
        .Q(n2573) );
  AO22X1 U2458 ( .IN1(n6790), .IN2(n6351), .IN3(\FIFO[62][27] ), .IN4(n6356), 
        .Q(n2574) );
  AO22X1 U2459 ( .IN1(n6779), .IN2(n6351), .IN3(\FIFO[62][28] ), .IN4(n6356), 
        .Q(n2575) );
  AO22X1 U2460 ( .IN1(n6768), .IN2(n6352), .IN3(\FIFO[62][29] ), .IN4(n6356), 
        .Q(n2576) );
  AO22X1 U2461 ( .IN1(n6757), .IN2(n6351), .IN3(\FIFO[62][30] ), .IN4(n6356), 
        .Q(n2577) );
  AO22X1 U2462 ( .IN1(n6746), .IN2(n6352), .IN3(\FIFO[62][31] ), .IN4(n6356), 
        .Q(n2578) );
  AO21X1 U2463 ( .IN1(n323), .IN2(n241), .IN3(n5973), .Q(n324) );
  AO22X1 U2464 ( .IN1(n7093), .IN2(n6347), .IN3(\FIFO[61][0] ), .IN4(n6348), 
        .Q(n2579) );
  AO22X1 U2465 ( .IN1(n7076), .IN2(n6347), .IN3(\FIFO[61][1] ), .IN4(n6348), 
        .Q(n2580) );
  AO22X1 U2466 ( .IN1(n7065), .IN2(n6347), .IN3(\FIFO[61][2] ), .IN4(n6348), 
        .Q(n2581) );
  AO22X1 U2467 ( .IN1(n7054), .IN2(n6347), .IN3(\FIFO[61][3] ), .IN4(n6348), 
        .Q(n2582) );
  AO22X1 U2468 ( .IN1(n7043), .IN2(n6347), .IN3(\FIFO[61][4] ), .IN4(n6348), 
        .Q(n2583) );
  AO22X1 U2469 ( .IN1(n7032), .IN2(n6347), .IN3(\FIFO[61][5] ), .IN4(n6348), 
        .Q(n2584) );
  AO22X1 U2470 ( .IN1(n7021), .IN2(n6347), .IN3(\FIFO[61][6] ), .IN4(n6348), 
        .Q(n2585) );
  AO22X1 U2471 ( .IN1(n7010), .IN2(n6346), .IN3(\FIFO[61][7] ), .IN4(n6348), 
        .Q(n2586) );
  AO22X1 U2472 ( .IN1(n6999), .IN2(n6346), .IN3(\FIFO[61][8] ), .IN4(n6348), 
        .Q(n2587) );
  AO22X1 U2473 ( .IN1(n6988), .IN2(n6346), .IN3(\FIFO[61][9] ), .IN4(n6348), 
        .Q(n2588) );
  AO22X1 U2474 ( .IN1(n6977), .IN2(n6346), .IN3(\FIFO[61][10] ), .IN4(n6348), 
        .Q(n2589) );
  AO22X1 U2475 ( .IN1(n6966), .IN2(n6346), .IN3(\FIFO[61][11] ), .IN4(n6348), 
        .Q(n2590) );
  AO22X1 U2476 ( .IN1(n6955), .IN2(n6346), .IN3(\FIFO[61][12] ), .IN4(n6349), 
        .Q(n2591) );
  AO22X1 U2477 ( .IN1(n6944), .IN2(n6346), .IN3(\FIFO[61][13] ), .IN4(n6349), 
        .Q(n2592) );
  AO22X1 U2478 ( .IN1(n6933), .IN2(n6345), .IN3(\FIFO[61][14] ), .IN4(n6349), 
        .Q(n2593) );
  AO22X1 U2479 ( .IN1(n6922), .IN2(n6345), .IN3(\FIFO[61][15] ), .IN4(n6349), 
        .Q(n2594) );
  AO22X1 U2480 ( .IN1(n6911), .IN2(n6345), .IN3(\FIFO[61][16] ), .IN4(n6349), 
        .Q(n2595) );
  AO22X1 U2481 ( .IN1(n6900), .IN2(n6345), .IN3(\FIFO[61][17] ), .IN4(n6349), 
        .Q(n2596) );
  AO22X1 U2482 ( .IN1(n6889), .IN2(n6345), .IN3(\FIFO[61][18] ), .IN4(n6349), 
        .Q(n2597) );
  AO22X1 U2483 ( .IN1(n6878), .IN2(n6345), .IN3(\FIFO[61][19] ), .IN4(n6349), 
        .Q(n2598) );
  AO22X1 U2484 ( .IN1(n6867), .IN2(n6345), .IN3(\FIFO[61][20] ), .IN4(n6349), 
        .Q(n2599) );
  AO22X1 U2485 ( .IN1(n6856), .IN2(n6347), .IN3(\FIFO[61][21] ), .IN4(n6349), 
        .Q(n2600) );
  AO22X1 U2486 ( .IN1(n6845), .IN2(n6346), .IN3(\FIFO[61][22] ), .IN4(n6349), 
        .Q(n2601) );
  AO22X1 U2487 ( .IN1(n6834), .IN2(n6345), .IN3(\FIFO[61][23] ), .IN4(n6349), 
        .Q(n2602) );
  AO22X1 U2488 ( .IN1(n6823), .IN2(n325), .IN3(\FIFO[61][24] ), .IN4(n6350), 
        .Q(n2603) );
  AO22X1 U2489 ( .IN1(n6812), .IN2(n325), .IN3(\FIFO[61][25] ), .IN4(n6350), 
        .Q(n2604) );
  AO22X1 U2490 ( .IN1(n6801), .IN2(n325), .IN3(\FIFO[61][26] ), .IN4(n6350), 
        .Q(n2605) );
  AO22X1 U2491 ( .IN1(n6790), .IN2(n6347), .IN3(\FIFO[61][27] ), .IN4(n6350), 
        .Q(n2606) );
  AO22X1 U2492 ( .IN1(n6779), .IN2(n6346), .IN3(\FIFO[61][28] ), .IN4(n6350), 
        .Q(n2607) );
  AO22X1 U2493 ( .IN1(n6768), .IN2(n6347), .IN3(\FIFO[61][29] ), .IN4(n6350), 
        .Q(n2608) );
  AO22X1 U2494 ( .IN1(n6757), .IN2(n6346), .IN3(\FIFO[61][30] ), .IN4(n6350), 
        .Q(n2609) );
  AO22X1 U2495 ( .IN1(n6746), .IN2(n6345), .IN3(\FIFO[61][31] ), .IN4(n6350), 
        .Q(n2610) );
  AO22X1 U2497 ( .IN1(n7093), .IN2(n6341), .IN3(\FIFO[60][0] ), .IN4(n6342), 
        .Q(n2611) );
  AO22X1 U2498 ( .IN1(n7076), .IN2(n6341), .IN3(\FIFO[60][1] ), .IN4(n6342), 
        .Q(n2612) );
  AO22X1 U2499 ( .IN1(n7065), .IN2(n6341), .IN3(\FIFO[60][2] ), .IN4(n6342), 
        .Q(n2613) );
  AO22X1 U2500 ( .IN1(n7054), .IN2(n6341), .IN3(\FIFO[60][3] ), .IN4(n6342), 
        .Q(n2614) );
  AO22X1 U2501 ( .IN1(n7043), .IN2(n6341), .IN3(\FIFO[60][4] ), .IN4(n6342), 
        .Q(n2615) );
  AO22X1 U2502 ( .IN1(n7032), .IN2(n6341), .IN3(\FIFO[60][5] ), .IN4(n6342), 
        .Q(n2616) );
  AO22X1 U2503 ( .IN1(n7021), .IN2(n6341), .IN3(\FIFO[60][6] ), .IN4(n6342), 
        .Q(n2617) );
  AO22X1 U2504 ( .IN1(n7010), .IN2(n6340), .IN3(\FIFO[60][7] ), .IN4(n6342), 
        .Q(n2618) );
  AO22X1 U2505 ( .IN1(n6999), .IN2(n6340), .IN3(\FIFO[60][8] ), .IN4(n6342), 
        .Q(n2619) );
  AO22X1 U2506 ( .IN1(n6988), .IN2(n6340), .IN3(\FIFO[60][9] ), .IN4(n6342), 
        .Q(n2620) );
  AO22X1 U2507 ( .IN1(n6977), .IN2(n6340), .IN3(\FIFO[60][10] ), .IN4(n6342), 
        .Q(n2621) );
  AO22X1 U2508 ( .IN1(n6966), .IN2(n6340), .IN3(\FIFO[60][11] ), .IN4(n6342), 
        .Q(n2622) );
  AO22X1 U2509 ( .IN1(n6955), .IN2(n6340), .IN3(\FIFO[60][12] ), .IN4(n6343), 
        .Q(n2623) );
  AO22X1 U2510 ( .IN1(n6944), .IN2(n6340), .IN3(\FIFO[60][13] ), .IN4(n6343), 
        .Q(n2624) );
  AO22X1 U2511 ( .IN1(n6933), .IN2(n6339), .IN3(\FIFO[60][14] ), .IN4(n6343), 
        .Q(n2625) );
  AO22X1 U2512 ( .IN1(n6922), .IN2(n6339), .IN3(\FIFO[60][15] ), .IN4(n6343), 
        .Q(n2626) );
  AO22X1 U2513 ( .IN1(n6911), .IN2(n6339), .IN3(\FIFO[60][16] ), .IN4(n6343), 
        .Q(n2627) );
  AO22X1 U2514 ( .IN1(n6900), .IN2(n6339), .IN3(\FIFO[60][17] ), .IN4(n6343), 
        .Q(n2628) );
  AO22X1 U2515 ( .IN1(n6889), .IN2(n6339), .IN3(\FIFO[60][18] ), .IN4(n6343), 
        .Q(n2629) );
  AO22X1 U2516 ( .IN1(n6878), .IN2(n6339), .IN3(\FIFO[60][19] ), .IN4(n6343), 
        .Q(n2630) );
  AO22X1 U2517 ( .IN1(n6867), .IN2(n6339), .IN3(\FIFO[60][20] ), .IN4(n6343), 
        .Q(n2631) );
  AO22X1 U2518 ( .IN1(n6856), .IN2(n6341), .IN3(\FIFO[60][21] ), .IN4(n6343), 
        .Q(n2632) );
  AO22X1 U2519 ( .IN1(n6845), .IN2(n6340), .IN3(\FIFO[60][22] ), .IN4(n6343), 
        .Q(n2633) );
  AO22X1 U2520 ( .IN1(n6834), .IN2(n6339), .IN3(\FIFO[60][23] ), .IN4(n6343), 
        .Q(n2634) );
  AO22X1 U2521 ( .IN1(n6823), .IN2(n326), .IN3(\FIFO[60][24] ), .IN4(n6344), 
        .Q(n2635) );
  AO22X1 U2522 ( .IN1(n6812), .IN2(n326), .IN3(\FIFO[60][25] ), .IN4(n6344), 
        .Q(n2636) );
  AO22X1 U2523 ( .IN1(n6801), .IN2(n326), .IN3(\FIFO[60][26] ), .IN4(n6344), 
        .Q(n2637) );
  AO22X1 U2524 ( .IN1(n6790), .IN2(n6341), .IN3(\FIFO[60][27] ), .IN4(n6344), 
        .Q(n2638) );
  AO22X1 U2525 ( .IN1(n6779), .IN2(n6340), .IN3(\FIFO[60][28] ), .IN4(n6344), 
        .Q(n2639) );
  AO22X1 U2526 ( .IN1(n6768), .IN2(n6341), .IN3(\FIFO[60][29] ), .IN4(n6344), 
        .Q(n2640) );
  AO22X1 U2527 ( .IN1(n6757), .IN2(n6340), .IN3(\FIFO[60][30] ), .IN4(n6344), 
        .Q(n2641) );
  AO22X1 U2528 ( .IN1(n6746), .IN2(n6339), .IN3(\FIFO[60][31] ), .IN4(n6344), 
        .Q(n2642) );
  AO21X1 U2529 ( .IN1(n323), .IN2(n245), .IN3(n7360), .Q(n326) );
  AO22X1 U2554 ( .IN1(n6822), .IN2(n327), .IN3(\FIFO[59][24] ), .IN4(n6338), 
        .Q(n2667) );
  AO22X1 U2555 ( .IN1(n6811), .IN2(n327), .IN3(\FIFO[59][25] ), .IN4(n6338), 
        .Q(n2668) );
  AO22X1 U2556 ( .IN1(n6800), .IN2(n327), .IN3(\FIFO[59][26] ), .IN4(n6338), 
        .Q(n2669) );
  AO22X1 U2557 ( .IN1(n6789), .IN2(n6335), .IN3(\FIFO[59][27] ), .IN4(n6338), 
        .Q(n2670) );
  AO22X1 U2558 ( .IN1(n6778), .IN2(n6335), .IN3(\FIFO[59][28] ), .IN4(n6338), 
        .Q(n2671) );
  AO22X1 U2559 ( .IN1(n6767), .IN2(n6334), .IN3(\FIFO[59][29] ), .IN4(n6338), 
        .Q(n2672) );
  AO22X1 U2560 ( .IN1(n6756), .IN2(n6333), .IN3(\FIFO[59][30] ), .IN4(n6338), 
        .Q(n2673) );
  AO22X1 U2561 ( .IN1(n6745), .IN2(n6334), .IN3(\FIFO[59][31] ), .IN4(n6338), 
        .Q(n2674) );
  AO21X1 U2562 ( .IN1(n323), .IN2(n247), .IN3(n7360), .Q(n327) );
  AO22X1 U2587 ( .IN1(n6822), .IN2(n6327), .IN3(\FIFO[58][24] ), .IN4(n6332), 
        .Q(n2699) );
  AO22X1 U2588 ( .IN1(n6811), .IN2(n6327), .IN3(\FIFO[58][25] ), .IN4(n6332), 
        .Q(n2700) );
  AO22X1 U2589 ( .IN1(n6800), .IN2(n6327), .IN3(\FIFO[58][26] ), .IN4(n6332), 
        .Q(n2701) );
  AO22X1 U2590 ( .IN1(n6789), .IN2(n6327), .IN3(\FIFO[58][27] ), .IN4(n6332), 
        .Q(n2702) );
  AO22X1 U2591 ( .IN1(n6778), .IN2(n6327), .IN3(\FIFO[58][28] ), .IN4(n6332), 
        .Q(n2703) );
  AO22X1 U2592 ( .IN1(n6767), .IN2(n6328), .IN3(\FIFO[58][29] ), .IN4(n6332), 
        .Q(n2704) );
  AO22X1 U2593 ( .IN1(n6756), .IN2(n6327), .IN3(\FIFO[58][30] ), .IN4(n6332), 
        .Q(n2705) );
  AO22X1 U2594 ( .IN1(n6745), .IN2(n6328), .IN3(\FIFO[58][31] ), .IN4(n6332), 
        .Q(n2706) );
  AO21X1 U2595 ( .IN1(n323), .IN2(n249), .IN3(n7360), .Q(n328) );
  AO22X1 U2596 ( .IN1(n7092), .IN2(n6323), .IN3(\FIFO[57][0] ), .IN4(n6324), 
        .Q(n2707) );
  AO22X1 U2597 ( .IN1(n7075), .IN2(n6322), .IN3(\FIFO[57][1] ), .IN4(n6324), 
        .Q(n2708) );
  AO22X1 U2599 ( .IN1(n7053), .IN2(n6323), .IN3(\FIFO[57][3] ), .IN4(n6324), 
        .Q(n2710) );
  AO22X1 U2600 ( .IN1(n7042), .IN2(n6322), .IN3(\FIFO[57][4] ), .IN4(n6324), 
        .Q(n2711) );
  AO22X1 U2601 ( .IN1(n7031), .IN2(n6321), .IN3(\FIFO[57][5] ), .IN4(n6324), 
        .Q(n2712) );
  AO22X1 U2602 ( .IN1(n7020), .IN2(n6323), .IN3(\FIFO[57][6] ), .IN4(n6324), 
        .Q(n2713) );
  AO22X1 U2603 ( .IN1(n7009), .IN2(n6323), .IN3(\FIFO[57][7] ), .IN4(n6324), 
        .Q(n2714) );
  AO22X1 U2604 ( .IN1(n6998), .IN2(n6323), .IN3(\FIFO[57][8] ), .IN4(n6324), 
        .Q(n2715) );
  AO22X1 U2605 ( .IN1(n6987), .IN2(n6323), .IN3(\FIFO[57][9] ), .IN4(n6324), 
        .Q(n2716) );
  AO22X1 U2606 ( .IN1(n6976), .IN2(n6323), .IN3(\FIFO[57][10] ), .IN4(n6324), 
        .Q(n2717) );
  AO22X1 U2607 ( .IN1(n6965), .IN2(n6323), .IN3(\FIFO[57][11] ), .IN4(n6324), 
        .Q(n2718) );
  AO22X1 U2608 ( .IN1(n6954), .IN2(n6323), .IN3(\FIFO[57][12] ), .IN4(n6325), 
        .Q(n2719) );
  AO22X1 U2609 ( .IN1(n6943), .IN2(n6323), .IN3(\FIFO[57][13] ), .IN4(n6325), 
        .Q(n2720) );
  AO22X1 U2610 ( .IN1(n6932), .IN2(n6322), .IN3(\FIFO[57][14] ), .IN4(n6325), 
        .Q(n2721) );
  AO22X1 U2611 ( .IN1(n6921), .IN2(n6322), .IN3(\FIFO[57][15] ), .IN4(n6325), 
        .Q(n2722) );
  AO22X1 U2612 ( .IN1(n6910), .IN2(n6322), .IN3(\FIFO[57][16] ), .IN4(n6325), 
        .Q(n2723) );
  AO22X1 U2614 ( .IN1(n6888), .IN2(n6322), .IN3(\FIFO[57][18] ), .IN4(n6325), 
        .Q(n2725) );
  AO22X1 U2615 ( .IN1(n6877), .IN2(n6322), .IN3(\FIFO[57][19] ), .IN4(n6325), 
        .Q(n2726) );
  AO22X1 U2616 ( .IN1(n6866), .IN2(n6322), .IN3(\FIFO[57][20] ), .IN4(n6325), 
        .Q(n2727) );
  AO22X1 U2617 ( .IN1(n6855), .IN2(n6321), .IN3(\FIFO[57][21] ), .IN4(n6325), 
        .Q(n2728) );
  AO22X1 U2618 ( .IN1(n6844), .IN2(n6321), .IN3(\FIFO[57][22] ), .IN4(n6325), 
        .Q(n2729) );
  AO22X1 U2619 ( .IN1(n6833), .IN2(n6321), .IN3(\FIFO[57][23] ), .IN4(n6325), 
        .Q(n2730) );
  AO22X1 U2620 ( .IN1(n6822), .IN2(n6321), .IN3(\FIFO[57][24] ), .IN4(n6326), 
        .Q(n2731) );
  AO22X1 U2621 ( .IN1(n6811), .IN2(n6321), .IN3(\FIFO[57][25] ), .IN4(n6326), 
        .Q(n2732) );
  AO22X1 U2622 ( .IN1(n6800), .IN2(n6321), .IN3(\FIFO[57][26] ), .IN4(n6326), 
        .Q(n2733) );
  AO22X1 U2623 ( .IN1(n6789), .IN2(n6321), .IN3(\FIFO[57][27] ), .IN4(n6326), 
        .Q(n2734) );
  AO22X1 U2624 ( .IN1(n6778), .IN2(n6321), .IN3(\FIFO[57][28] ), .IN4(n6326), 
        .Q(n2735) );
  AO22X1 U2625 ( .IN1(n6767), .IN2(n6322), .IN3(\FIFO[57][29] ), .IN4(n6326), 
        .Q(n2736) );
  AO22X1 U2626 ( .IN1(n6756), .IN2(n6321), .IN3(\FIFO[57][30] ), .IN4(n6326), 
        .Q(n2737) );
  AO22X1 U2627 ( .IN1(n6745), .IN2(n6322), .IN3(\FIFO[57][31] ), .IN4(n6326), 
        .Q(n2738) );
  AO21X1 U2628 ( .IN1(n323), .IN2(n251), .IN3(n7360), .Q(n329) );
  AO22X1 U2629 ( .IN1(n7092), .IN2(n6317), .IN3(\FIFO[56][0] ), .IN4(n6318), 
        .Q(n2739) );
  AO22X1 U2630 ( .IN1(n7075), .IN2(n6317), .IN3(\FIFO[56][1] ), .IN4(n6318), 
        .Q(n2740) );
  AO22X1 U2631 ( .IN1(n7064), .IN2(n6317), .IN3(\FIFO[56][2] ), .IN4(n6318), 
        .Q(n2741) );
  AO22X1 U2632 ( .IN1(n7053), .IN2(n6317), .IN3(\FIFO[56][3] ), .IN4(n6318), 
        .Q(n2742) );
  AO22X1 U2633 ( .IN1(n7042), .IN2(n6317), .IN3(\FIFO[56][4] ), .IN4(n6318), 
        .Q(n2743) );
  AO22X1 U2634 ( .IN1(n7031), .IN2(n6317), .IN3(\FIFO[56][5] ), .IN4(n6318), 
        .Q(n2744) );
  AO22X1 U2635 ( .IN1(n7020), .IN2(n6317), .IN3(\FIFO[56][6] ), .IN4(n6318), 
        .Q(n2745) );
  AO22X1 U2636 ( .IN1(n7009), .IN2(n6316), .IN3(\FIFO[56][7] ), .IN4(n6318), 
        .Q(n2746) );
  AO22X1 U2637 ( .IN1(n6998), .IN2(n6316), .IN3(\FIFO[56][8] ), .IN4(n6318), 
        .Q(n2747) );
  AO22X1 U2638 ( .IN1(n6987), .IN2(n6316), .IN3(\FIFO[56][9] ), .IN4(n6318), 
        .Q(n2748) );
  AO22X1 U2639 ( .IN1(n6976), .IN2(n6316), .IN3(\FIFO[56][10] ), .IN4(n6318), 
        .Q(n2749) );
  AO22X1 U2640 ( .IN1(n6965), .IN2(n6316), .IN3(\FIFO[56][11] ), .IN4(n6318), 
        .Q(n2750) );
  AO22X1 U2641 ( .IN1(n6954), .IN2(n6316), .IN3(\FIFO[56][12] ), .IN4(n6319), 
        .Q(n2751) );
  AO22X1 U2642 ( .IN1(n6943), .IN2(n6316), .IN3(\FIFO[56][13] ), .IN4(n6319), 
        .Q(n2752) );
  AO22X1 U2643 ( .IN1(n6932), .IN2(n6315), .IN3(\FIFO[56][14] ), .IN4(n6319), 
        .Q(n2753) );
  AO22X1 U2644 ( .IN1(n6921), .IN2(n6315), .IN3(\FIFO[56][15] ), .IN4(n6319), 
        .Q(n2754) );
  AO22X1 U2645 ( .IN1(n6910), .IN2(n6315), .IN3(\FIFO[56][16] ), .IN4(n6319), 
        .Q(n2755) );
  AO22X1 U2646 ( .IN1(n6899), .IN2(n6315), .IN3(\FIFO[56][17] ), .IN4(n6319), 
        .Q(n2756) );
  AO22X1 U2647 ( .IN1(n6888), .IN2(n6315), .IN3(\FIFO[56][18] ), .IN4(n6319), 
        .Q(n2757) );
  AO22X1 U2648 ( .IN1(n6877), .IN2(n6315), .IN3(\FIFO[56][19] ), .IN4(n6319), 
        .Q(n2758) );
  AO22X1 U2649 ( .IN1(n6866), .IN2(n6315), .IN3(\FIFO[56][20] ), .IN4(n6319), 
        .Q(n2759) );
  AO22X1 U2650 ( .IN1(n6855), .IN2(n6317), .IN3(\FIFO[56][21] ), .IN4(n6319), 
        .Q(n2760) );
  AO22X1 U2651 ( .IN1(n6844), .IN2(n6316), .IN3(\FIFO[56][22] ), .IN4(n6319), 
        .Q(n2761) );
  AO22X1 U2652 ( .IN1(n6833), .IN2(n6315), .IN3(\FIFO[56][23] ), .IN4(n6319), 
        .Q(n2762) );
  AO22X1 U2653 ( .IN1(n6822), .IN2(n330), .IN3(\FIFO[56][24] ), .IN4(n6320), 
        .Q(n2763) );
  AO22X1 U2654 ( .IN1(n6811), .IN2(n330), .IN3(\FIFO[56][25] ), .IN4(n6320), 
        .Q(n2764) );
  AO22X1 U2655 ( .IN1(n6800), .IN2(n330), .IN3(\FIFO[56][26] ), .IN4(n6320), 
        .Q(n2765) );
  AO22X1 U2656 ( .IN1(n6789), .IN2(n6317), .IN3(\FIFO[56][27] ), .IN4(n6320), 
        .Q(n2766) );
  AO22X1 U2657 ( .IN1(n6778), .IN2(n6316), .IN3(\FIFO[56][28] ), .IN4(n6320), 
        .Q(n2767) );
  AO22X1 U2658 ( .IN1(n6767), .IN2(n6317), .IN3(\FIFO[56][29] ), .IN4(n6320), 
        .Q(n2768) );
  AO22X1 U2659 ( .IN1(n6756), .IN2(n6316), .IN3(\FIFO[56][30] ), .IN4(n6320), 
        .Q(n2769) );
  AO22X1 U2660 ( .IN1(n6745), .IN2(n6315), .IN3(\FIFO[56][31] ), .IN4(n6320), 
        .Q(n2770) );
  AO21X1 U2661 ( .IN1(n323), .IN2(n253), .IN3(n7360), .Q(n330) );
  AO22X1 U2686 ( .IN1(n6822), .IN2(n331), .IN3(\FIFO[55][24] ), .IN4(n6314), 
        .Q(n2795) );
  AO22X1 U2687 ( .IN1(n6811), .IN2(n331), .IN3(\FIFO[55][25] ), .IN4(n6314), 
        .Q(n2796) );
  AO22X1 U2688 ( .IN1(n6800), .IN2(n331), .IN3(\FIFO[55][26] ), .IN4(n6314), 
        .Q(n2797) );
  AO22X1 U2689 ( .IN1(n6789), .IN2(n6311), .IN3(\FIFO[55][27] ), .IN4(n6314), 
        .Q(n2798) );
  AO22X1 U2690 ( .IN1(n6778), .IN2(n6310), .IN3(\FIFO[55][28] ), .IN4(n6314), 
        .Q(n2799) );
  AO22X1 U2691 ( .IN1(n6767), .IN2(n6311), .IN3(\FIFO[55][29] ), .IN4(n6314), 
        .Q(n2800) );
  AO22X1 U2692 ( .IN1(n6756), .IN2(n6310), .IN3(\FIFO[55][30] ), .IN4(n6314), 
        .Q(n2801) );
  AO22X1 U2693 ( .IN1(n6745), .IN2(n6309), .IN3(\FIFO[55][31] ), .IN4(n6314), 
        .Q(n2802) );
  AO21X1 U2694 ( .IN1(n323), .IN2(n255), .IN3(n7360), .Q(n331) );
  AO22X1 U2719 ( .IN1(n6822), .IN2(n332), .IN3(\FIFO[54][24] ), .IN4(n6308), 
        .Q(n2827) );
  AO22X1 U2720 ( .IN1(n6811), .IN2(n332), .IN3(\FIFO[54][25] ), .IN4(n6308), 
        .Q(n2828) );
  AO22X1 U2721 ( .IN1(n6800), .IN2(n332), .IN3(\FIFO[54][26] ), .IN4(n6308), 
        .Q(n2829) );
  AO22X1 U2722 ( .IN1(n6789), .IN2(n6305), .IN3(\FIFO[54][27] ), .IN4(n6308), 
        .Q(n2830) );
  AO22X1 U2723 ( .IN1(n6778), .IN2(n6305), .IN3(\FIFO[54][28] ), .IN4(n6308), 
        .Q(n2831) );
  AO22X1 U2724 ( .IN1(n6767), .IN2(n6304), .IN3(\FIFO[54][29] ), .IN4(n6308), 
        .Q(n2832) );
  AO22X1 U2725 ( .IN1(n6756), .IN2(n6303), .IN3(\FIFO[54][30] ), .IN4(n6308), 
        .Q(n2833) );
  AO22X1 U2726 ( .IN1(n6745), .IN2(n6304), .IN3(\FIFO[54][31] ), .IN4(n6308), 
        .Q(n2834) );
  AO21X1 U2727 ( .IN1(n323), .IN2(n257), .IN3(n7360), .Q(n332) );
  AO22X1 U2728 ( .IN1(n7092), .IN2(n6299), .IN3(\FIFO[53][0] ), .IN4(n6300), 
        .Q(n2835) );
  AO22X1 U2729 ( .IN1(n7075), .IN2(n6299), .IN3(\FIFO[53][1] ), .IN4(n6300), 
        .Q(n2836) );
  AO22X1 U2730 ( .IN1(n7064), .IN2(n6299), .IN3(\FIFO[53][2] ), .IN4(n6300), 
        .Q(n2837) );
  AO22X1 U2731 ( .IN1(n7053), .IN2(n6299), .IN3(\FIFO[53][3] ), .IN4(n6300), 
        .Q(n2838) );
  AO22X1 U2732 ( .IN1(n7042), .IN2(n6299), .IN3(\FIFO[53][4] ), .IN4(n6300), 
        .Q(n2839) );
  AO22X1 U2733 ( .IN1(n7031), .IN2(n6299), .IN3(\FIFO[53][5] ), .IN4(n6300), 
        .Q(n2840) );
  AO22X1 U2734 ( .IN1(n7020), .IN2(n6299), .IN3(\FIFO[53][6] ), .IN4(n6300), 
        .Q(n2841) );
  AO22X1 U2735 ( .IN1(n7009), .IN2(n6298), .IN3(\FIFO[53][7] ), .IN4(n6300), 
        .Q(n2842) );
  AO22X1 U2736 ( .IN1(n6998), .IN2(n6298), .IN3(\FIFO[53][8] ), .IN4(n6300), 
        .Q(n2843) );
  AO22X1 U2737 ( .IN1(n6987), .IN2(n6298), .IN3(\FIFO[53][9] ), .IN4(n6300), 
        .Q(n2844) );
  AO22X1 U2738 ( .IN1(n6976), .IN2(n6298), .IN3(\FIFO[53][10] ), .IN4(n6300), 
        .Q(n2845) );
  AO22X1 U2739 ( .IN1(n6965), .IN2(n6298), .IN3(\FIFO[53][11] ), .IN4(n6300), 
        .Q(n2846) );
  AO22X1 U2740 ( .IN1(n6954), .IN2(n6298), .IN3(\FIFO[53][12] ), .IN4(n6301), 
        .Q(n2847) );
  AO22X1 U2741 ( .IN1(n6943), .IN2(n6298), .IN3(\FIFO[53][13] ), .IN4(n6301), 
        .Q(n2848) );
  AO22X1 U2742 ( .IN1(n6932), .IN2(n6299), .IN3(\FIFO[53][14] ), .IN4(n6301), 
        .Q(n2849) );
  AO22X1 U2743 ( .IN1(n6921), .IN2(n6298), .IN3(\FIFO[53][15] ), .IN4(n6301), 
        .Q(n2850) );
  AO22X1 U2744 ( .IN1(n6910), .IN2(n6297), .IN3(\FIFO[53][16] ), .IN4(n6301), 
        .Q(n2851) );
  AO22X1 U2745 ( .IN1(n6899), .IN2(n6299), .IN3(\FIFO[53][17] ), .IN4(n6301), 
        .Q(n2852) );
  AO22X1 U2747 ( .IN1(n6877), .IN2(n6297), .IN3(\FIFO[53][19] ), .IN4(n6301), 
        .Q(n2854) );
  AO22X1 U2748 ( .IN1(n6866), .IN2(n6299), .IN3(\FIFO[53][20] ), .IN4(n6301), 
        .Q(n2855) );
  AO22X1 U2749 ( .IN1(n6855), .IN2(n6297), .IN3(\FIFO[53][21] ), .IN4(n6301), 
        .Q(n2856) );
  AO22X1 U2750 ( .IN1(n6844), .IN2(n6297), .IN3(\FIFO[53][22] ), .IN4(n6301), 
        .Q(n2857) );
  AO22X1 U2751 ( .IN1(n6833), .IN2(n6297), .IN3(\FIFO[53][23] ), .IN4(n6301), 
        .Q(n2858) );
  AO22X1 U2752 ( .IN1(n6822), .IN2(n6297), .IN3(\FIFO[53][24] ), .IN4(n6302), 
        .Q(n2859) );
  AO22X1 U2753 ( .IN1(n6811), .IN2(n6297), .IN3(\FIFO[53][25] ), .IN4(n6302), 
        .Q(n2860) );
  AO22X1 U2754 ( .IN1(n6800), .IN2(n6297), .IN3(\FIFO[53][26] ), .IN4(n6302), 
        .Q(n2861) );
  AO22X1 U2755 ( .IN1(n6789), .IN2(n6297), .IN3(\FIFO[53][27] ), .IN4(n6302), 
        .Q(n2862) );
  AO22X1 U2756 ( .IN1(n6778), .IN2(n6297), .IN3(\FIFO[53][28] ), .IN4(n6302), 
        .Q(n2863) );
  AO22X1 U2757 ( .IN1(n6767), .IN2(n6298), .IN3(\FIFO[53][29] ), .IN4(n6302), 
        .Q(n2864) );
  AO22X1 U2758 ( .IN1(n6756), .IN2(n6297), .IN3(\FIFO[53][30] ), .IN4(n6302), 
        .Q(n2865) );
  AO22X1 U2759 ( .IN1(n6745), .IN2(n6298), .IN3(\FIFO[53][31] ), .IN4(n6302), 
        .Q(n2866) );
  AO21X1 U2760 ( .IN1(n323), .IN2(n259), .IN3(n7360), .Q(n333) );
  AO22X1 U2761 ( .IN1(n7092), .IN2(n6293), .IN3(\FIFO[52][0] ), .IN4(n6294), 
        .Q(n2867) );
  AO22X1 U2762 ( .IN1(n7075), .IN2(n6292), .IN3(\FIFO[52][1] ), .IN4(n6294), 
        .Q(n2868) );
  AO22X1 U2763 ( .IN1(n7064), .IN2(n6291), .IN3(\FIFO[52][2] ), .IN4(n6294), 
        .Q(n2869) );
  AO22X1 U2764 ( .IN1(n7053), .IN2(n6293), .IN3(\FIFO[52][3] ), .IN4(n6294), 
        .Q(n2870) );
  AO22X1 U2765 ( .IN1(n7042), .IN2(n6292), .IN3(\FIFO[52][4] ), .IN4(n6294), 
        .Q(n2871) );
  AO22X1 U2767 ( .IN1(n7020), .IN2(n6293), .IN3(\FIFO[52][6] ), .IN4(n6294), 
        .Q(n2873) );
  AO22X1 U2768 ( .IN1(n7009), .IN2(n6293), .IN3(\FIFO[52][7] ), .IN4(n6294), 
        .Q(n2874) );
  AO22X1 U2769 ( .IN1(n6998), .IN2(n6293), .IN3(\FIFO[52][8] ), .IN4(n6294), 
        .Q(n2875) );
  AO22X1 U2770 ( .IN1(n6987), .IN2(n6293), .IN3(\FIFO[52][9] ), .IN4(n6294), 
        .Q(n2876) );
  AO22X1 U2771 ( .IN1(n6976), .IN2(n6293), .IN3(\FIFO[52][10] ), .IN4(n6294), 
        .Q(n2877) );
  AO22X1 U2772 ( .IN1(n6965), .IN2(n6293), .IN3(\FIFO[52][11] ), .IN4(n6294), 
        .Q(n2878) );
  AO22X1 U2773 ( .IN1(n6954), .IN2(n6293), .IN3(\FIFO[52][12] ), .IN4(n6295), 
        .Q(n2879) );
  AO22X1 U2774 ( .IN1(n6943), .IN2(n6293), .IN3(\FIFO[52][13] ), .IN4(n6295), 
        .Q(n2880) );
  AO22X1 U2775 ( .IN1(n6932), .IN2(n6292), .IN3(\FIFO[52][14] ), .IN4(n6295), 
        .Q(n2881) );
  AO22X1 U2776 ( .IN1(n6921), .IN2(n6292), .IN3(\FIFO[52][15] ), .IN4(n6295), 
        .Q(n2882) );
  AO22X1 U2777 ( .IN1(n6910), .IN2(n6292), .IN3(\FIFO[52][16] ), .IN4(n6295), 
        .Q(n2883) );
  AO22X1 U2778 ( .IN1(n6899), .IN2(n6292), .IN3(\FIFO[52][17] ), .IN4(n6295), 
        .Q(n2884) );
  AO22X1 U2779 ( .IN1(n6888), .IN2(n6292), .IN3(\FIFO[52][18] ), .IN4(n6295), 
        .Q(n2885) );
  AO22X1 U2781 ( .IN1(n6866), .IN2(n6292), .IN3(\FIFO[52][20] ), .IN4(n6295), 
        .Q(n2887) );
  AO22X1 U2782 ( .IN1(n6855), .IN2(n6291), .IN3(\FIFO[52][21] ), .IN4(n6295), 
        .Q(n2888) );
  AO22X1 U2783 ( .IN1(n6844), .IN2(n6291), .IN3(\FIFO[52][22] ), .IN4(n6295), 
        .Q(n2889) );
  AO22X1 U2784 ( .IN1(n6833), .IN2(n6291), .IN3(\FIFO[52][23] ), .IN4(n6295), 
        .Q(n2890) );
  AO22X1 U2785 ( .IN1(n6822), .IN2(n6291), .IN3(\FIFO[52][24] ), .IN4(n6296), 
        .Q(n2891) );
  AO22X1 U2786 ( .IN1(n6811), .IN2(n6291), .IN3(\FIFO[52][25] ), .IN4(n6296), 
        .Q(n2892) );
  AO22X1 U2787 ( .IN1(n6800), .IN2(n6291), .IN3(\FIFO[52][26] ), .IN4(n6296), 
        .Q(n2893) );
  AO22X1 U2788 ( .IN1(n6789), .IN2(n6291), .IN3(\FIFO[52][27] ), .IN4(n6296), 
        .Q(n2894) );
  AO22X1 U2789 ( .IN1(n6778), .IN2(n6291), .IN3(\FIFO[52][28] ), .IN4(n6296), 
        .Q(n2895) );
  AO22X1 U2790 ( .IN1(n6767), .IN2(n6292), .IN3(\FIFO[52][29] ), .IN4(n6296), 
        .Q(n2896) );
  AO22X1 U2791 ( .IN1(n6756), .IN2(n6291), .IN3(\FIFO[52][30] ), .IN4(n6296), 
        .Q(n2897) );
  AO22X1 U2792 ( .IN1(n6745), .IN2(n6292), .IN3(\FIFO[52][31] ), .IN4(n6296), 
        .Q(n2898) );
  AO21X1 U2793 ( .IN1(n323), .IN2(n261), .IN3(n7360), .Q(n334) );
  AO22X1 U2818 ( .IN1(n6822), .IN2(n335), .IN3(\FIFO[51][24] ), .IN4(n6290), 
        .Q(n2923) );
  AO22X1 U2819 ( .IN1(n6811), .IN2(n335), .IN3(\FIFO[51][25] ), .IN4(n6290), 
        .Q(n2924) );
  AO22X1 U2820 ( .IN1(n6800), .IN2(n335), .IN3(\FIFO[51][26] ), .IN4(n6290), 
        .Q(n2925) );
  AO22X1 U2821 ( .IN1(n6789), .IN2(n6287), .IN3(\FIFO[51][27] ), .IN4(n6290), 
        .Q(n2926) );
  AO22X1 U2822 ( .IN1(n6778), .IN2(n6286), .IN3(\FIFO[51][28] ), .IN4(n6290), 
        .Q(n2927) );
  AO22X1 U2823 ( .IN1(n6767), .IN2(n6287), .IN3(\FIFO[51][29] ), .IN4(n6290), 
        .Q(n2928) );
  AO22X1 U2824 ( .IN1(n6756), .IN2(n6286), .IN3(\FIFO[51][30] ), .IN4(n6290), 
        .Q(n2929) );
  AO22X1 U2825 ( .IN1(n6745), .IN2(n6285), .IN3(\FIFO[51][31] ), .IN4(n6290), 
        .Q(n2930) );
  AO21X1 U2826 ( .IN1(n323), .IN2(n263), .IN3(n7360), .Q(n335) );
  AO22X1 U2851 ( .IN1(n6822), .IN2(n336), .IN3(\FIFO[50][24] ), .IN4(n6284), 
        .Q(n2955) );
  AO22X1 U2852 ( .IN1(n6811), .IN2(n336), .IN3(\FIFO[50][25] ), .IN4(n6284), 
        .Q(n2956) );
  AO22X1 U2853 ( .IN1(n6800), .IN2(n336), .IN3(\FIFO[50][26] ), .IN4(n6284), 
        .Q(n2957) );
  AO22X1 U2854 ( .IN1(n6789), .IN2(n6281), .IN3(\FIFO[50][27] ), .IN4(n6284), 
        .Q(n2958) );
  AO22X1 U2855 ( .IN1(n6778), .IN2(n6280), .IN3(\FIFO[50][28] ), .IN4(n6284), 
        .Q(n2959) );
  AO22X1 U2856 ( .IN1(n6767), .IN2(n6281), .IN3(\FIFO[50][29] ), .IN4(n6284), 
        .Q(n2960) );
  AO22X1 U2857 ( .IN1(n6756), .IN2(n6280), .IN3(\FIFO[50][30] ), .IN4(n6284), 
        .Q(n2961) );
  AO22X1 U2858 ( .IN1(n6745), .IN2(n6279), .IN3(\FIFO[50][31] ), .IN4(n6284), 
        .Q(n2962) );
  AO21X1 U2859 ( .IN1(n323), .IN2(n265), .IN3(n7360), .Q(n336) );
  AO22X1 U2860 ( .IN1(n7092), .IN2(n6275), .IN3(\FIFO[49][0] ), .IN4(n6276), 
        .Q(n2963) );
  AO22X1 U2861 ( .IN1(n7075), .IN2(n6275), .IN3(\FIFO[49][1] ), .IN4(n6276), 
        .Q(n2964) );
  AO22X1 U2862 ( .IN1(n7064), .IN2(n6275), .IN3(\FIFO[49][2] ), .IN4(n6276), 
        .Q(n2965) );
  AO22X1 U2863 ( .IN1(n7053), .IN2(n6275), .IN3(\FIFO[49][3] ), .IN4(n6276), 
        .Q(n2966) );
  AO22X1 U2864 ( .IN1(n7042), .IN2(n6275), .IN3(\FIFO[49][4] ), .IN4(n6276), 
        .Q(n2967) );
  AO22X1 U2865 ( .IN1(n7031), .IN2(n6275), .IN3(\FIFO[49][5] ), .IN4(n6276), 
        .Q(n2968) );
  AO22X1 U2866 ( .IN1(n7020), .IN2(n6275), .IN3(\FIFO[49][6] ), .IN4(n6276), 
        .Q(n2969) );
  AO22X1 U2867 ( .IN1(n7009), .IN2(n6274), .IN3(\FIFO[49][7] ), .IN4(n6276), 
        .Q(n2970) );
  AO22X1 U2868 ( .IN1(n6998), .IN2(n6274), .IN3(\FIFO[49][8] ), .IN4(n6276), 
        .Q(n2971) );
  AO22X1 U2869 ( .IN1(n6987), .IN2(n6274), .IN3(\FIFO[49][9] ), .IN4(n6276), 
        .Q(n2972) );
  AO22X1 U2870 ( .IN1(n6976), .IN2(n6274), .IN3(\FIFO[49][10] ), .IN4(n6276), 
        .Q(n2973) );
  AO22X1 U2871 ( .IN1(n6965), .IN2(n6274), .IN3(\FIFO[49][11] ), .IN4(n6276), 
        .Q(n2974) );
  AO22X1 U2872 ( .IN1(n6954), .IN2(n6274), .IN3(\FIFO[49][12] ), .IN4(n6277), 
        .Q(n2975) );
  AO22X1 U2873 ( .IN1(n6943), .IN2(n6274), .IN3(\FIFO[49][13] ), .IN4(n6277), 
        .Q(n2976) );
  AO22X1 U2874 ( .IN1(n6932), .IN2(n6273), .IN3(\FIFO[49][14] ), .IN4(n6277), 
        .Q(n2977) );
  AO22X1 U2875 ( .IN1(n6921), .IN2(n6273), .IN3(\FIFO[49][15] ), .IN4(n6277), 
        .Q(n2978) );
  AO22X1 U2876 ( .IN1(n6910), .IN2(n6273), .IN3(\FIFO[49][16] ), .IN4(n6277), 
        .Q(n2979) );
  AO22X1 U2877 ( .IN1(n6899), .IN2(n6273), .IN3(\FIFO[49][17] ), .IN4(n6277), 
        .Q(n2980) );
  AO22X1 U2878 ( .IN1(n6888), .IN2(n6273), .IN3(\FIFO[49][18] ), .IN4(n6277), 
        .Q(n2981) );
  AO22X1 U2879 ( .IN1(n6877), .IN2(n6273), .IN3(\FIFO[49][19] ), .IN4(n6277), 
        .Q(n2982) );
  AO22X1 U2880 ( .IN1(n6866), .IN2(n6273), .IN3(\FIFO[49][20] ), .IN4(n6277), 
        .Q(n2983) );
  AO22X1 U2881 ( .IN1(n6855), .IN2(n6275), .IN3(\FIFO[49][21] ), .IN4(n6277), 
        .Q(n2984) );
  AO22X1 U2882 ( .IN1(n6844), .IN2(n6274), .IN3(\FIFO[49][22] ), .IN4(n6277), 
        .Q(n2985) );
  AO22X1 U2883 ( .IN1(n6833), .IN2(n6273), .IN3(\FIFO[49][23] ), .IN4(n6277), 
        .Q(n2986) );
  AO22X1 U2884 ( .IN1(n6822), .IN2(n337), .IN3(\FIFO[49][24] ), .IN4(n6278), 
        .Q(n2987) );
  AO22X1 U2885 ( .IN1(n6811), .IN2(n337), .IN3(\FIFO[49][25] ), .IN4(n6278), 
        .Q(n2988) );
  AO22X1 U2886 ( .IN1(n6800), .IN2(n337), .IN3(\FIFO[49][26] ), .IN4(n6278), 
        .Q(n2989) );
  AO22X1 U2887 ( .IN1(n6789), .IN2(n6275), .IN3(\FIFO[49][27] ), .IN4(n6278), 
        .Q(n2990) );
  AO22X1 U2888 ( .IN1(n6778), .IN2(n6275), .IN3(\FIFO[49][28] ), .IN4(n6278), 
        .Q(n2991) );
  AO22X1 U2889 ( .IN1(n6767), .IN2(n6274), .IN3(\FIFO[49][29] ), .IN4(n6278), 
        .Q(n2992) );
  AO22X1 U2890 ( .IN1(n6756), .IN2(n6273), .IN3(\FIFO[49][30] ), .IN4(n6278), 
        .Q(n2993) );
  AO22X1 U2891 ( .IN1(n6745), .IN2(n6274), .IN3(\FIFO[49][31] ), .IN4(n6278), 
        .Q(n2994) );
  AO21X1 U2892 ( .IN1(n323), .IN2(n267), .IN3(n7360), .Q(n337) );
  AO22X1 U2893 ( .IN1(n7092), .IN2(n6269), .IN3(\FIFO[48][0] ), .IN4(n6270), 
        .Q(n2995) );
  AO22X1 U2894 ( .IN1(n7075), .IN2(n6269), .IN3(\FIFO[48][1] ), .IN4(n6270), 
        .Q(n2996) );
  AO22X1 U2895 ( .IN1(n7064), .IN2(n6269), .IN3(\FIFO[48][2] ), .IN4(n6270), 
        .Q(n2997) );
  AO22X1 U2896 ( .IN1(n7053), .IN2(n6269), .IN3(\FIFO[48][3] ), .IN4(n6270), 
        .Q(n2998) );
  AO22X1 U2897 ( .IN1(n7042), .IN2(n6269), .IN3(\FIFO[48][4] ), .IN4(n6270), 
        .Q(n2999) );
  AO22X1 U2898 ( .IN1(n7031), .IN2(n6269), .IN3(\FIFO[48][5] ), .IN4(n6270), 
        .Q(n3000) );
  AO22X1 U2899 ( .IN1(n7020), .IN2(n6269), .IN3(\FIFO[48][6] ), .IN4(n6270), 
        .Q(n3001) );
  AO22X1 U2900 ( .IN1(n7009), .IN2(n6268), .IN3(\FIFO[48][7] ), .IN4(n6270), 
        .Q(n3002) );
  AO22X1 U2901 ( .IN1(n6998), .IN2(n6268), .IN3(\FIFO[48][8] ), .IN4(n6270), 
        .Q(n3003) );
  AO22X1 U2902 ( .IN1(n6987), .IN2(n6268), .IN3(\FIFO[48][9] ), .IN4(n6270), 
        .Q(n3004) );
  AO22X1 U2903 ( .IN1(n6976), .IN2(n6268), .IN3(\FIFO[48][10] ), .IN4(n6270), 
        .Q(n3005) );
  AO22X1 U2905 ( .IN1(n6954), .IN2(n6268), .IN3(\FIFO[48][12] ), .IN4(n6271), 
        .Q(n3007) );
  AO22X1 U2906 ( .IN1(n6943), .IN2(n6268), .IN3(\FIFO[48][13] ), .IN4(n6271), 
        .Q(n3008) );
  AO22X1 U2907 ( .IN1(n6932), .IN2(n6269), .IN3(\FIFO[48][14] ), .IN4(n6271), 
        .Q(n3009) );
  AO22X1 U2908 ( .IN1(n6921), .IN2(n6268), .IN3(\FIFO[48][15] ), .IN4(n6271), 
        .Q(n3010) );
  AO22X1 U2909 ( .IN1(n6910), .IN2(n6267), .IN3(\FIFO[48][16] ), .IN4(n6271), 
        .Q(n3011) );
  AO22X1 U2910 ( .IN1(n6899), .IN2(n6269), .IN3(\FIFO[48][17] ), .IN4(n6271), 
        .Q(n3012) );
  AO22X1 U2911 ( .IN1(n6888), .IN2(n6268), .IN3(\FIFO[48][18] ), .IN4(n6271), 
        .Q(n3013) );
  AO22X1 U2912 ( .IN1(n6877), .IN2(n6267), .IN3(\FIFO[48][19] ), .IN4(n6271), 
        .Q(n3014) );
  AO22X1 U2914 ( .IN1(n6855), .IN2(n6267), .IN3(\FIFO[48][21] ), .IN4(n6271), 
        .Q(n3016) );
  AO22X1 U2915 ( .IN1(n6844), .IN2(n6267), .IN3(\FIFO[48][22] ), .IN4(n6271), 
        .Q(n3017) );
  AO22X1 U2916 ( .IN1(n6833), .IN2(n6267), .IN3(\FIFO[48][23] ), .IN4(n6271), 
        .Q(n3018) );
  AO22X1 U2917 ( .IN1(n6822), .IN2(n6267), .IN3(\FIFO[48][24] ), .IN4(n6272), 
        .Q(n3019) );
  AO22X1 U2918 ( .IN1(n6811), .IN2(n6267), .IN3(\FIFO[48][25] ), .IN4(n6272), 
        .Q(n3020) );
  AO22X1 U2919 ( .IN1(n6800), .IN2(n6267), .IN3(\FIFO[48][26] ), .IN4(n6272), 
        .Q(n3021) );
  AO22X1 U2920 ( .IN1(n6789), .IN2(n6267), .IN3(\FIFO[48][27] ), .IN4(n6272), 
        .Q(n3022) );
  AO22X1 U2921 ( .IN1(n6778), .IN2(n6267), .IN3(\FIFO[48][28] ), .IN4(n6272), 
        .Q(n3023) );
  AO22X1 U2922 ( .IN1(n6767), .IN2(n6268), .IN3(\FIFO[48][29] ), .IN4(n6272), 
        .Q(n3024) );
  AO22X1 U2923 ( .IN1(n6756), .IN2(n6267), .IN3(\FIFO[48][30] ), .IN4(n6272), 
        .Q(n3025) );
  AO22X1 U2924 ( .IN1(n6745), .IN2(n6268), .IN3(\FIFO[48][31] ), .IN4(n6272), 
        .Q(n3026) );
  AO21X1 U2925 ( .IN1(n323), .IN2(n269), .IN3(n7360), .Q(n338) );
  AO22X1 U2951 ( .IN1(n6821), .IN2(n339), .IN3(\FIFO[47][24] ), .IN4(n6266), 
        .Q(n3051) );
  AO22X1 U2952 ( .IN1(n6810), .IN2(n339), .IN3(\FIFO[47][25] ), .IN4(n6266), 
        .Q(n3052) );
  AO22X1 U2953 ( .IN1(n6799), .IN2(n339), .IN3(\FIFO[47][26] ), .IN4(n6266), 
        .Q(n3053) );
  AO22X1 U2954 ( .IN1(n6788), .IN2(n6263), .IN3(\FIFO[47][27] ), .IN4(n6266), 
        .Q(n3054) );
  AO22X1 U2955 ( .IN1(n6777), .IN2(n6262), .IN3(\FIFO[47][28] ), .IN4(n6266), 
        .Q(n3055) );
  AO22X1 U2956 ( .IN1(n6766), .IN2(n6263), .IN3(\FIFO[47][29] ), .IN4(n6266), 
        .Q(n3056) );
  AO22X1 U2957 ( .IN1(n6755), .IN2(n6262), .IN3(\FIFO[47][30] ), .IN4(n6266), 
        .Q(n3057) );
  AO22X1 U2958 ( .IN1(n6744), .IN2(n6261), .IN3(\FIFO[47][31] ), .IN4(n6266), 
        .Q(n3058) );
  AO21X1 U2959 ( .IN1(n340), .IN2(n238), .IN3(n7360), .Q(n339) );
  AO22X1 U2984 ( .IN1(n6821), .IN2(n341), .IN3(\FIFO[46][24] ), .IN4(n6260), 
        .Q(n3083) );
  AO22X1 U2985 ( .IN1(n6810), .IN2(n341), .IN3(\FIFO[46][25] ), .IN4(n6260), 
        .Q(n3084) );
  AO22X1 U2986 ( .IN1(n6799), .IN2(n341), .IN3(\FIFO[46][26] ), .IN4(n6260), 
        .Q(n3085) );
  AO22X1 U2987 ( .IN1(n6788), .IN2(n6257), .IN3(\FIFO[46][27] ), .IN4(n6260), 
        .Q(n3086) );
  AO22X1 U2988 ( .IN1(n6777), .IN2(n6256), .IN3(\FIFO[46][28] ), .IN4(n6260), 
        .Q(n3087) );
  AO22X1 U2989 ( .IN1(n6766), .IN2(n6257), .IN3(\FIFO[46][29] ), .IN4(n6260), 
        .Q(n3088) );
  AO22X1 U2990 ( .IN1(n6755), .IN2(n6256), .IN3(\FIFO[46][30] ), .IN4(n6260), 
        .Q(n3089) );
  AO22X1 U2991 ( .IN1(n6744), .IN2(n6255), .IN3(\FIFO[46][31] ), .IN4(n6260), 
        .Q(n3090) );
  AO21X1 U2992 ( .IN1(n340), .IN2(n241), .IN3(n7360), .Q(n341) );
  AO22X1 U2993 ( .IN1(n7091), .IN2(n6251), .IN3(\FIFO[45][0] ), .IN4(n6252), 
        .Q(n3091) );
  AO22X1 U2994 ( .IN1(n7074), .IN2(n6251), .IN3(\FIFO[45][1] ), .IN4(n6252), 
        .Q(n3092) );
  AO22X1 U2995 ( .IN1(n7063), .IN2(n6251), .IN3(\FIFO[45][2] ), .IN4(n6252), 
        .Q(n3093) );
  AO22X1 U2996 ( .IN1(n7052), .IN2(n6251), .IN3(\FIFO[45][3] ), .IN4(n6252), 
        .Q(n3094) );
  AO22X1 U2997 ( .IN1(n7041), .IN2(n6251), .IN3(\FIFO[45][4] ), .IN4(n6252), 
        .Q(n3095) );
  AO22X1 U2998 ( .IN1(n7030), .IN2(n6251), .IN3(\FIFO[45][5] ), .IN4(n6252), 
        .Q(n3096) );
  AO22X1 U2999 ( .IN1(n7019), .IN2(n6251), .IN3(\FIFO[45][6] ), .IN4(n6252), 
        .Q(n3097) );
  AO22X1 U3000 ( .IN1(n7008), .IN2(n6250), .IN3(\FIFO[45][7] ), .IN4(n6252), 
        .Q(n3098) );
  AO22X1 U3001 ( .IN1(n6997), .IN2(n6250), .IN3(\FIFO[45][8] ), .IN4(n6252), 
        .Q(n3099) );
  AO22X1 U3002 ( .IN1(n6986), .IN2(n6250), .IN3(\FIFO[45][9] ), .IN4(n6252), 
        .Q(n3100) );
  AO22X1 U3003 ( .IN1(n6975), .IN2(n6250), .IN3(\FIFO[45][10] ), .IN4(n6252), 
        .Q(n3101) );
  AO22X1 U3004 ( .IN1(n6964), .IN2(n6250), .IN3(\FIFO[45][11] ), .IN4(n6252), 
        .Q(n3102) );
  AO22X1 U3005 ( .IN1(n6953), .IN2(n6250), .IN3(\FIFO[45][12] ), .IN4(n6253), 
        .Q(n3103) );
  AO22X1 U3006 ( .IN1(n6942), .IN2(n6250), .IN3(\FIFO[45][13] ), .IN4(n6253), 
        .Q(n3104) );
  AO22X1 U3007 ( .IN1(n6931), .IN2(n6249), .IN3(\FIFO[45][14] ), .IN4(n6253), 
        .Q(n3105) );
  AO22X1 U3008 ( .IN1(n6920), .IN2(n6249), .IN3(\FIFO[45][15] ), .IN4(n6253), 
        .Q(n3106) );
  AO22X1 U3009 ( .IN1(n6909), .IN2(n6249), .IN3(\FIFO[45][16] ), .IN4(n6253), 
        .Q(n3107) );
  AO22X1 U3010 ( .IN1(n6898), .IN2(n6249), .IN3(\FIFO[45][17] ), .IN4(n6253), 
        .Q(n3108) );
  AO22X1 U3011 ( .IN1(n6887), .IN2(n6249), .IN3(\FIFO[45][18] ), .IN4(n6253), 
        .Q(n3109) );
  AO22X1 U3012 ( .IN1(n6876), .IN2(n6249), .IN3(\FIFO[45][19] ), .IN4(n6253), 
        .Q(n3110) );
  AO22X1 U3013 ( .IN1(n6865), .IN2(n6249), .IN3(\FIFO[45][20] ), .IN4(n6253), 
        .Q(n3111) );
  AO22X1 U3014 ( .IN1(n6854), .IN2(n6251), .IN3(\FIFO[45][21] ), .IN4(n6253), 
        .Q(n3112) );
  AO22X1 U3015 ( .IN1(n6843), .IN2(n6250), .IN3(\FIFO[45][22] ), .IN4(n6253), 
        .Q(n3113) );
  AO22X1 U3016 ( .IN1(n6832), .IN2(n6249), .IN3(\FIFO[45][23] ), .IN4(n6253), 
        .Q(n3114) );
  AO22X1 U3017 ( .IN1(n6821), .IN2(n342), .IN3(\FIFO[45][24] ), .IN4(n6254), 
        .Q(n3115) );
  AO22X1 U3018 ( .IN1(n6810), .IN2(n342), .IN3(\FIFO[45][25] ), .IN4(n6254), 
        .Q(n3116) );
  AO22X1 U3019 ( .IN1(n6799), .IN2(n342), .IN3(\FIFO[45][26] ), .IN4(n6254), 
        .Q(n3117) );
  AO22X1 U3020 ( .IN1(n6788), .IN2(n6251), .IN3(\FIFO[45][27] ), .IN4(n6254), 
        .Q(n3118) );
  AO22X1 U3021 ( .IN1(n6777), .IN2(n6251), .IN3(\FIFO[45][28] ), .IN4(n6254), 
        .Q(n3119) );
  AO22X1 U3022 ( .IN1(n6766), .IN2(n6250), .IN3(\FIFO[45][29] ), .IN4(n6254), 
        .Q(n3120) );
  AO22X1 U3023 ( .IN1(n6755), .IN2(n6249), .IN3(\FIFO[45][30] ), .IN4(n6254), 
        .Q(n3121) );
  AO22X1 U3024 ( .IN1(n6744), .IN2(n6250), .IN3(\FIFO[45][31] ), .IN4(n6254), 
        .Q(n3122) );
  AO21X1 U3025 ( .IN1(n340), .IN2(n243), .IN3(n7360), .Q(n342) );
  AO22X1 U3027 ( .IN1(n7074), .IN2(n6245), .IN3(\FIFO[44][1] ), .IN4(n6246), 
        .Q(n3124) );
  AO22X1 U3028 ( .IN1(n7063), .IN2(n6245), .IN3(\FIFO[44][2] ), .IN4(n6246), 
        .Q(n3125) );
  AO22X1 U3029 ( .IN1(n7052), .IN2(n6245), .IN3(\FIFO[44][3] ), .IN4(n6246), 
        .Q(n3126) );
  AO22X1 U3030 ( .IN1(n7041), .IN2(n6245), .IN3(\FIFO[44][4] ), .IN4(n6246), 
        .Q(n3127) );
  AO22X1 U3031 ( .IN1(n7030), .IN2(n6245), .IN3(\FIFO[44][5] ), .IN4(n6246), 
        .Q(n3128) );
  AO22X1 U3032 ( .IN1(n7019), .IN2(n6245), .IN3(\FIFO[44][6] ), .IN4(n6246), 
        .Q(n3129) );
  AO22X1 U3033 ( .IN1(n7008), .IN2(n6244), .IN3(\FIFO[44][7] ), .IN4(n6246), 
        .Q(n3130) );
  AO22X1 U3034 ( .IN1(n6997), .IN2(n6244), .IN3(\FIFO[44][8] ), .IN4(n6246), 
        .Q(n3131) );
  AO22X1 U3035 ( .IN1(n6986), .IN2(n6244), .IN3(\FIFO[44][9] ), .IN4(n6246), 
        .Q(n3132) );
  AO22X1 U3036 ( .IN1(n6975), .IN2(n6244), .IN3(\FIFO[44][10] ), .IN4(n6246), 
        .Q(n3133) );
  AO22X1 U3037 ( .IN1(n6964), .IN2(n6244), .IN3(\FIFO[44][11] ), .IN4(n6246), 
        .Q(n3134) );
  AO22X1 U3038 ( .IN1(n6953), .IN2(n6244), .IN3(\FIFO[44][12] ), .IN4(n6247), 
        .Q(n3135) );
  AO22X1 U3039 ( .IN1(n6942), .IN2(n6244), .IN3(\FIFO[44][13] ), .IN4(n6247), 
        .Q(n3136) );
  AO22X1 U3040 ( .IN1(n6931), .IN2(n6245), .IN3(\FIFO[44][14] ), .IN4(n6247), 
        .Q(n3137) );
  AO22X1 U3041 ( .IN1(n6920), .IN2(n6244), .IN3(\FIFO[44][15] ), .IN4(n6247), 
        .Q(n3138) );
  AO22X1 U3042 ( .IN1(n6909), .IN2(n6243), .IN3(\FIFO[44][16] ), .IN4(n6247), 
        .Q(n3139) );
  AO22X1 U3043 ( .IN1(n6898), .IN2(n6245), .IN3(\FIFO[44][17] ), .IN4(n6247), 
        .Q(n3140) );
  AO22X1 U3044 ( .IN1(n6887), .IN2(n6244), .IN3(\FIFO[44][18] ), .IN4(n6247), 
        .Q(n3141) );
  AO22X1 U3045 ( .IN1(n6876), .IN2(n6243), .IN3(\FIFO[44][19] ), .IN4(n6247), 
        .Q(n3142) );
  AO22X1 U3046 ( .IN1(n6865), .IN2(n6245), .IN3(\FIFO[44][20] ), .IN4(n6247), 
        .Q(n3143) );
  AO22X1 U3048 ( .IN1(n6843), .IN2(n6243), .IN3(\FIFO[44][22] ), .IN4(n6247), 
        .Q(n3145) );
  AO22X1 U3049 ( .IN1(n6832), .IN2(n6243), .IN3(\FIFO[44][23] ), .IN4(n6247), 
        .Q(n3146) );
  AO22X1 U3050 ( .IN1(n6821), .IN2(n6243), .IN3(\FIFO[44][24] ), .IN4(n6248), 
        .Q(n3147) );
  AO22X1 U3051 ( .IN1(n6810), .IN2(n6243), .IN3(\FIFO[44][25] ), .IN4(n6248), 
        .Q(n3148) );
  AO22X1 U3052 ( .IN1(n6799), .IN2(n6243), .IN3(\FIFO[44][26] ), .IN4(n6248), 
        .Q(n3149) );
  AO22X1 U3053 ( .IN1(n6788), .IN2(n6243), .IN3(\FIFO[44][27] ), .IN4(n6248), 
        .Q(n3150) );
  AO22X1 U3054 ( .IN1(n6777), .IN2(n6243), .IN3(\FIFO[44][28] ), .IN4(n6248), 
        .Q(n3151) );
  AO22X1 U3055 ( .IN1(n6766), .IN2(n6244), .IN3(\FIFO[44][29] ), .IN4(n6248), 
        .Q(n3152) );
  AO22X1 U3056 ( .IN1(n6755), .IN2(n6243), .IN3(\FIFO[44][30] ), .IN4(n6248), 
        .Q(n3153) );
  AO22X1 U3057 ( .IN1(n6744), .IN2(n6244), .IN3(\FIFO[44][31] ), .IN4(n6248), 
        .Q(n3154) );
  AO21X1 U3058 ( .IN1(n340), .IN2(n245), .IN3(n7360), .Q(n343) );
  AO22X1 U3083 ( .IN1(n6821), .IN2(n6237), .IN3(\FIFO[43][24] ), .IN4(n6242), 
        .Q(n3179) );
  AO22X1 U3084 ( .IN1(n6810), .IN2(n6237), .IN3(\FIFO[43][25] ), .IN4(n6242), 
        .Q(n3180) );
  AO22X1 U3085 ( .IN1(n6799), .IN2(n6237), .IN3(\FIFO[43][26] ), .IN4(n6242), 
        .Q(n3181) );
  AO22X1 U3086 ( .IN1(n6788), .IN2(n6237), .IN3(\FIFO[43][27] ), .IN4(n6242), 
        .Q(n3182) );
  AO22X1 U3087 ( .IN1(n6777), .IN2(n6237), .IN3(\FIFO[43][28] ), .IN4(n6242), 
        .Q(n3183) );
  AO22X1 U3088 ( .IN1(n6766), .IN2(n6238), .IN3(\FIFO[43][29] ), .IN4(n6242), 
        .Q(n3184) );
  AO22X1 U3089 ( .IN1(n6755), .IN2(n6237), .IN3(\FIFO[43][30] ), .IN4(n6242), 
        .Q(n3185) );
  AO22X1 U3090 ( .IN1(n6744), .IN2(n6238), .IN3(\FIFO[43][31] ), .IN4(n6242), 
        .Q(n3186) );
  AO21X1 U3091 ( .IN1(n340), .IN2(n247), .IN3(n7360), .Q(n344) );
  AO22X1 U3116 ( .IN1(n6821), .IN2(n345), .IN3(\FIFO[42][24] ), .IN4(n6236), 
        .Q(n3211) );
  AO22X1 U3117 ( .IN1(n6810), .IN2(n345), .IN3(\FIFO[42][25] ), .IN4(n6236), 
        .Q(n3212) );
  AO22X1 U3118 ( .IN1(n6799), .IN2(n345), .IN3(\FIFO[42][26] ), .IN4(n6236), 
        .Q(n3213) );
  AO22X1 U3119 ( .IN1(n6788), .IN2(n6233), .IN3(\FIFO[42][27] ), .IN4(n6236), 
        .Q(n3214) );
  AO22X1 U3120 ( .IN1(n6777), .IN2(n6232), .IN3(\FIFO[42][28] ), .IN4(n6236), 
        .Q(n3215) );
  AO22X1 U3121 ( .IN1(n6766), .IN2(n6233), .IN3(\FIFO[42][29] ), .IN4(n6236), 
        .Q(n3216) );
  AO22X1 U3122 ( .IN1(n6755), .IN2(n6232), .IN3(\FIFO[42][30] ), .IN4(n6236), 
        .Q(n3217) );
  AO22X1 U3123 ( .IN1(n6744), .IN2(n6231), .IN3(\FIFO[42][31] ), .IN4(n6236), 
        .Q(n3218) );
  AO21X1 U3124 ( .IN1(n340), .IN2(n249), .IN3(n7360), .Q(n345) );
  AO22X1 U3125 ( .IN1(n7091), .IN2(n6227), .IN3(\FIFO[41][0] ), .IN4(n6228), 
        .Q(n3219) );
  AO22X1 U3126 ( .IN1(n7074), .IN2(n6227), .IN3(\FIFO[41][1] ), .IN4(n6228), 
        .Q(n3220) );
  AO22X1 U3127 ( .IN1(n7063), .IN2(n6227), .IN3(\FIFO[41][2] ), .IN4(n6228), 
        .Q(n3221) );
  AO22X1 U3128 ( .IN1(n7052), .IN2(n6227), .IN3(\FIFO[41][3] ), .IN4(n6228), 
        .Q(n3222) );
  AO22X1 U3129 ( .IN1(n7041), .IN2(n6227), .IN3(\FIFO[41][4] ), .IN4(n6228), 
        .Q(n3223) );
  AO22X1 U3130 ( .IN1(n7030), .IN2(n6227), .IN3(\FIFO[41][5] ), .IN4(n6228), 
        .Q(n3224) );
  AO22X1 U3131 ( .IN1(n7019), .IN2(n6227), .IN3(\FIFO[41][6] ), .IN4(n6228), 
        .Q(n3225) );
  AO22X1 U3132 ( .IN1(n7008), .IN2(n6226), .IN3(\FIFO[41][7] ), .IN4(n6228), 
        .Q(n3226) );
  AO22X1 U3134 ( .IN1(n6986), .IN2(n6226), .IN3(\FIFO[41][9] ), .IN4(n6228), 
        .Q(n3228) );
  AO22X1 U3135 ( .IN1(n6975), .IN2(n6226), .IN3(\FIFO[41][10] ), .IN4(n6228), 
        .Q(n3229) );
  AO22X1 U3136 ( .IN1(n6964), .IN2(n6226), .IN3(\FIFO[41][11] ), .IN4(n6228), 
        .Q(n3230) );
  AO22X1 U3137 ( .IN1(n6953), .IN2(n6226), .IN3(\FIFO[41][12] ), .IN4(n6229), 
        .Q(n3231) );
  AO22X1 U3138 ( .IN1(n6942), .IN2(n6226), .IN3(\FIFO[41][13] ), .IN4(n6229), 
        .Q(n3232) );
  AO22X1 U3139 ( .IN1(n6931), .IN2(n6225), .IN3(\FIFO[41][14] ), .IN4(n6229), 
        .Q(n3233) );
  AO22X1 U3140 ( .IN1(n6920), .IN2(n6225), .IN3(\FIFO[41][15] ), .IN4(n6229), 
        .Q(n3234) );
  AO22X1 U3141 ( .IN1(n6909), .IN2(n6225), .IN3(\FIFO[41][16] ), .IN4(n6229), 
        .Q(n3235) );
  AO22X1 U3142 ( .IN1(n6898), .IN2(n6225), .IN3(\FIFO[41][17] ), .IN4(n6229), 
        .Q(n3236) );
  AO22X1 U3143 ( .IN1(n6887), .IN2(n6225), .IN3(\FIFO[41][18] ), .IN4(n6229), 
        .Q(n3237) );
  AO22X1 U3144 ( .IN1(n6876), .IN2(n6225), .IN3(\FIFO[41][19] ), .IN4(n6229), 
        .Q(n3238) );
  AO22X1 U3145 ( .IN1(n6865), .IN2(n6225), .IN3(\FIFO[41][20] ), .IN4(n6229), 
        .Q(n3239) );
  AO22X1 U3146 ( .IN1(n6854), .IN2(n6227), .IN3(\FIFO[41][21] ), .IN4(n6229), 
        .Q(n3240) );
  AO22X1 U3147 ( .IN1(n6843), .IN2(n6226), .IN3(\FIFO[41][22] ), .IN4(n6229), 
        .Q(n3241) );
  AO22X1 U3148 ( .IN1(n6832), .IN2(n6225), .IN3(\FIFO[41][23] ), .IN4(n6229), 
        .Q(n3242) );
  AO22X1 U3149 ( .IN1(n6821), .IN2(n346), .IN3(\FIFO[41][24] ), .IN4(n6230), 
        .Q(n3243) );
  AO22X1 U3150 ( .IN1(n6810), .IN2(n346), .IN3(\FIFO[41][25] ), .IN4(n6230), 
        .Q(n3244) );
  AO22X1 U3151 ( .IN1(n6799), .IN2(n346), .IN3(\FIFO[41][26] ), .IN4(n6230), 
        .Q(n3245) );
  AO22X1 U3152 ( .IN1(n6788), .IN2(n6227), .IN3(\FIFO[41][27] ), .IN4(n6230), 
        .Q(n3246) );
  AO22X1 U3153 ( .IN1(n6777), .IN2(n6226), .IN3(\FIFO[41][28] ), .IN4(n6230), 
        .Q(n3247) );
  AO22X1 U3154 ( .IN1(n6766), .IN2(n6227), .IN3(\FIFO[41][29] ), .IN4(n6230), 
        .Q(n3248) );
  AO22X1 U3155 ( .IN1(n6755), .IN2(n6226), .IN3(\FIFO[41][30] ), .IN4(n6230), 
        .Q(n3249) );
  AO22X1 U3156 ( .IN1(n6744), .IN2(n6225), .IN3(\FIFO[41][31] ), .IN4(n6230), 
        .Q(n3250) );
  AO21X1 U3157 ( .IN1(n340), .IN2(n251), .IN3(n7360), .Q(n346) );
  AO22X1 U3158 ( .IN1(n7091), .IN2(n6221), .IN3(\FIFO[40][0] ), .IN4(n6222), 
        .Q(n3251) );
  AO22X1 U3159 ( .IN1(n7074), .IN2(n6221), .IN3(\FIFO[40][1] ), .IN4(n6222), 
        .Q(n3252) );
  AO22X1 U3160 ( .IN1(n7063), .IN2(n6221), .IN3(\FIFO[40][2] ), .IN4(n6222), 
        .Q(n3253) );
  AO22X1 U3161 ( .IN1(n7052), .IN2(n6221), .IN3(\FIFO[40][3] ), .IN4(n6222), 
        .Q(n3254) );
  AO22X1 U3162 ( .IN1(n7041), .IN2(n6221), .IN3(\FIFO[40][4] ), .IN4(n6222), 
        .Q(n3255) );
  AO22X1 U3163 ( .IN1(n7030), .IN2(n6221), .IN3(\FIFO[40][5] ), .IN4(n6222), 
        .Q(n3256) );
  AO22X1 U3164 ( .IN1(n7019), .IN2(n6221), .IN3(\FIFO[40][6] ), .IN4(n6222), 
        .Q(n3257) );
  AO22X1 U3165 ( .IN1(n7008), .IN2(n6220), .IN3(\FIFO[40][7] ), .IN4(n6222), 
        .Q(n3258) );
  AO22X1 U3166 ( .IN1(n6997), .IN2(n6220), .IN3(\FIFO[40][8] ), .IN4(n6222), 
        .Q(n3259) );
  AO22X1 U3168 ( .IN1(n6975), .IN2(n6220), .IN3(\FIFO[40][10] ), .IN4(n6222), 
        .Q(n3261) );
  AO22X1 U3169 ( .IN1(n6964), .IN2(n6220), .IN3(\FIFO[40][11] ), .IN4(n6222), 
        .Q(n3262) );
  AO22X1 U3170 ( .IN1(n6953), .IN2(n6220), .IN3(\FIFO[40][12] ), .IN4(n6223), 
        .Q(n3263) );
  AO22X1 U3171 ( .IN1(n6942), .IN2(n6220), .IN3(\FIFO[40][13] ), .IN4(n6223), 
        .Q(n3264) );
  AO22X1 U3172 ( .IN1(n6931), .IN2(n6219), .IN3(\FIFO[40][14] ), .IN4(n6223), 
        .Q(n3265) );
  AO22X1 U3173 ( .IN1(n6920), .IN2(n6219), .IN3(\FIFO[40][15] ), .IN4(n6223), 
        .Q(n3266) );
  AO22X1 U3174 ( .IN1(n6909), .IN2(n6219), .IN3(\FIFO[40][16] ), .IN4(n6223), 
        .Q(n3267) );
  AO22X1 U3175 ( .IN1(n6898), .IN2(n6219), .IN3(\FIFO[40][17] ), .IN4(n6223), 
        .Q(n3268) );
  AO22X1 U3176 ( .IN1(n6887), .IN2(n6219), .IN3(\FIFO[40][18] ), .IN4(n6223), 
        .Q(n3269) );
  AO22X1 U3177 ( .IN1(n6876), .IN2(n6219), .IN3(\FIFO[40][19] ), .IN4(n6223), 
        .Q(n3270) );
  AO22X1 U3178 ( .IN1(n6865), .IN2(n6219), .IN3(\FIFO[40][20] ), .IN4(n6223), 
        .Q(n3271) );
  AO22X1 U3179 ( .IN1(n6854), .IN2(n6221), .IN3(\FIFO[40][21] ), .IN4(n6223), 
        .Q(n3272) );
  AO22X1 U3180 ( .IN1(n6843), .IN2(n6220), .IN3(\FIFO[40][22] ), .IN4(n6223), 
        .Q(n3273) );
  AO22X1 U3181 ( .IN1(n6832), .IN2(n6219), .IN3(\FIFO[40][23] ), .IN4(n6223), 
        .Q(n3274) );
  AO22X1 U3182 ( .IN1(n6821), .IN2(n347), .IN3(\FIFO[40][24] ), .IN4(n6224), 
        .Q(n3275) );
  AO22X1 U3183 ( .IN1(n6810), .IN2(n347), .IN3(\FIFO[40][25] ), .IN4(n6224), 
        .Q(n3276) );
  AO22X1 U3184 ( .IN1(n6799), .IN2(n347), .IN3(\FIFO[40][26] ), .IN4(n6224), 
        .Q(n3277) );
  AO22X1 U3185 ( .IN1(n6788), .IN2(n6221), .IN3(\FIFO[40][27] ), .IN4(n6224), 
        .Q(n3278) );
  AO22X1 U3186 ( .IN1(n6777), .IN2(n6221), .IN3(\FIFO[40][28] ), .IN4(n6224), 
        .Q(n3279) );
  AO22X1 U3187 ( .IN1(n6766), .IN2(n6220), .IN3(\FIFO[40][29] ), .IN4(n6224), 
        .Q(n3280) );
  AO22X1 U3188 ( .IN1(n6755), .IN2(n6219), .IN3(\FIFO[40][30] ), .IN4(n6224), 
        .Q(n3281) );
  AO22X1 U3189 ( .IN1(n6744), .IN2(n6220), .IN3(\FIFO[40][31] ), .IN4(n6224), 
        .Q(n3282) );
  AO21X1 U3190 ( .IN1(n340), .IN2(n253), .IN3(n7360), .Q(n347) );
  AO22X1 U3215 ( .IN1(n6821), .IN2(n6213), .IN3(\FIFO[39][24] ), .IN4(n6218), 
        .Q(n3307) );
  AO22X1 U3216 ( .IN1(n6810), .IN2(n6213), .IN3(\FIFO[39][25] ), .IN4(n6218), 
        .Q(n3308) );
  AO22X1 U3217 ( .IN1(n6799), .IN2(n6213), .IN3(\FIFO[39][26] ), .IN4(n6218), 
        .Q(n3309) );
  AO22X1 U3218 ( .IN1(n6788), .IN2(n6213), .IN3(\FIFO[39][27] ), .IN4(n6218), 
        .Q(n3310) );
  AO22X1 U3219 ( .IN1(n6777), .IN2(n6213), .IN3(\FIFO[39][28] ), .IN4(n6218), 
        .Q(n3311) );
  AO22X1 U3220 ( .IN1(n6766), .IN2(n6214), .IN3(\FIFO[39][29] ), .IN4(n6218), 
        .Q(n3312) );
  AO22X1 U3221 ( .IN1(n6755), .IN2(n6213), .IN3(\FIFO[39][30] ), .IN4(n6218), 
        .Q(n3313) );
  AO22X1 U3222 ( .IN1(n6744), .IN2(n6214), .IN3(\FIFO[39][31] ), .IN4(n6218), 
        .Q(n3314) );
  AO21X1 U3223 ( .IN1(n340), .IN2(n255), .IN3(n7360), .Q(n348) );
  AO22X1 U3249 ( .IN1(n6810), .IN2(n6207), .IN3(\FIFO[38][25] ), .IN4(n6212), 
        .Q(n3340) );
  AO22X1 U3250 ( .IN1(n6799), .IN2(n6207), .IN3(\FIFO[38][26] ), .IN4(n6212), 
        .Q(n3341) );
  AO22X1 U3251 ( .IN1(n6788), .IN2(n6207), .IN3(\FIFO[38][27] ), .IN4(n6212), 
        .Q(n3342) );
  AO22X1 U3252 ( .IN1(n6777), .IN2(n6207), .IN3(\FIFO[38][28] ), .IN4(n6212), 
        .Q(n3343) );
  AO22X1 U3253 ( .IN1(n6766), .IN2(n6208), .IN3(\FIFO[38][29] ), .IN4(n6212), 
        .Q(n3344) );
  AO22X1 U3254 ( .IN1(n6755), .IN2(n6207), .IN3(\FIFO[38][30] ), .IN4(n6212), 
        .Q(n3345) );
  AO22X1 U3255 ( .IN1(n6744), .IN2(n6208), .IN3(\FIFO[38][31] ), .IN4(n6212), 
        .Q(n3346) );
  AO21X1 U3256 ( .IN1(n340), .IN2(n257), .IN3(n7360), .Q(n349) );
  AO22X1 U3257 ( .IN1(n7091), .IN2(n6203), .IN3(\FIFO[37][0] ), .IN4(n6204), 
        .Q(n3347) );
  AO22X1 U3258 ( .IN1(n7074), .IN2(n6203), .IN3(\FIFO[37][1] ), .IN4(n6204), 
        .Q(n3348) );
  AO22X1 U3259 ( .IN1(n7063), .IN2(n6203), .IN3(\FIFO[37][2] ), .IN4(n6204), 
        .Q(n3349) );
  AO22X1 U3260 ( .IN1(n7052), .IN2(n6203), .IN3(\FIFO[37][3] ), .IN4(n6204), 
        .Q(n3350) );
  AO22X1 U3261 ( .IN1(n7041), .IN2(n6203), .IN3(\FIFO[37][4] ), .IN4(n6204), 
        .Q(n3351) );
  AO22X1 U3262 ( .IN1(n7030), .IN2(n6203), .IN3(\FIFO[37][5] ), .IN4(n6204), 
        .Q(n3352) );
  AO22X1 U3263 ( .IN1(n7019), .IN2(n6203), .IN3(\FIFO[37][6] ), .IN4(n6204), 
        .Q(n3353) );
  AO22X1 U3264 ( .IN1(n7008), .IN2(n6202), .IN3(\FIFO[37][7] ), .IN4(n6204), 
        .Q(n3354) );
  AO22X1 U3265 ( .IN1(n6997), .IN2(n6202), .IN3(\FIFO[37][8] ), .IN4(n6204), 
        .Q(n3355) );
  AO22X1 U3266 ( .IN1(n6986), .IN2(n6202), .IN3(\FIFO[37][9] ), .IN4(n6204), 
        .Q(n3356) );
  AO22X1 U3268 ( .IN1(n6964), .IN2(n6202), .IN3(\FIFO[37][11] ), .IN4(n6204), 
        .Q(n3358) );
  AO22X1 U3269 ( .IN1(n6953), .IN2(n6202), .IN3(\FIFO[37][12] ), .IN4(n6205), 
        .Q(n3359) );
  AO22X1 U3270 ( .IN1(n6942), .IN2(n6202), .IN3(\FIFO[37][13] ), .IN4(n6205), 
        .Q(n3360) );
  AO22X1 U3271 ( .IN1(n6931), .IN2(n6201), .IN3(\FIFO[37][14] ), .IN4(n6205), 
        .Q(n3361) );
  AO22X1 U3272 ( .IN1(n6920), .IN2(n6201), .IN3(\FIFO[37][15] ), .IN4(n6205), 
        .Q(n3362) );
  AO22X1 U3273 ( .IN1(n6909), .IN2(n6201), .IN3(\FIFO[37][16] ), .IN4(n6205), 
        .Q(n3363) );
  AO22X1 U3274 ( .IN1(n6898), .IN2(n6201), .IN3(\FIFO[37][17] ), .IN4(n6205), 
        .Q(n3364) );
  AO22X1 U3275 ( .IN1(n6887), .IN2(n6201), .IN3(\FIFO[37][18] ), .IN4(n6205), 
        .Q(n3365) );
  AO22X1 U3276 ( .IN1(n6876), .IN2(n6201), .IN3(\FIFO[37][19] ), .IN4(n6205), 
        .Q(n3366) );
  AO22X1 U3277 ( .IN1(n6865), .IN2(n6201), .IN3(\FIFO[37][20] ), .IN4(n6205), 
        .Q(n3367) );
  AO22X1 U3278 ( .IN1(n6854), .IN2(n6203), .IN3(\FIFO[37][21] ), .IN4(n6205), 
        .Q(n3368) );
  AO22X1 U3279 ( .IN1(n6843), .IN2(n6202), .IN3(\FIFO[37][22] ), .IN4(n6205), 
        .Q(n3369) );
  AO22X1 U3280 ( .IN1(n6832), .IN2(n6201), .IN3(\FIFO[37][23] ), .IN4(n6205), 
        .Q(n3370) );
  AO22X1 U3281 ( .IN1(n6821), .IN2(n350), .IN3(\FIFO[37][24] ), .IN4(n6206), 
        .Q(n3371) );
  AO22X1 U3282 ( .IN1(n6810), .IN2(n350), .IN3(\FIFO[37][25] ), .IN4(n6206), 
        .Q(n3372) );
  AO22X1 U3283 ( .IN1(n6799), .IN2(n350), .IN3(\FIFO[37][26] ), .IN4(n6206), 
        .Q(n3373) );
  AO22X1 U3284 ( .IN1(n6788), .IN2(n6203), .IN3(\FIFO[37][27] ), .IN4(n6206), 
        .Q(n3374) );
  AO22X1 U3285 ( .IN1(n6777), .IN2(n6202), .IN3(\FIFO[37][28] ), .IN4(n6206), 
        .Q(n3375) );
  AO22X1 U3286 ( .IN1(n6766), .IN2(n6203), .IN3(\FIFO[37][29] ), .IN4(n6206), 
        .Q(n3376) );
  AO22X1 U3287 ( .IN1(n6755), .IN2(n6202), .IN3(\FIFO[37][30] ), .IN4(n6206), 
        .Q(n3377) );
  AO22X1 U3288 ( .IN1(n6744), .IN2(n6201), .IN3(\FIFO[37][31] ), .IN4(n6206), 
        .Q(n3378) );
  AO21X1 U3289 ( .IN1(n340), .IN2(n259), .IN3(n7360), .Q(n350) );
  AO22X1 U3290 ( .IN1(n7091), .IN2(n6197), .IN3(\FIFO[36][0] ), .IN4(n6198), 
        .Q(n3379) );
  AO22X1 U3291 ( .IN1(n7074), .IN2(n6197), .IN3(\FIFO[36][1] ), .IN4(n6198), 
        .Q(n3380) );
  AO22X1 U3292 ( .IN1(n7063), .IN2(n6197), .IN3(\FIFO[36][2] ), .IN4(n6198), 
        .Q(n3381) );
  AO22X1 U3293 ( .IN1(n7052), .IN2(n6197), .IN3(\FIFO[36][3] ), .IN4(n6198), 
        .Q(n3382) );
  AO22X1 U3294 ( .IN1(n7041), .IN2(n6197), .IN3(\FIFO[36][4] ), .IN4(n6198), 
        .Q(n3383) );
  AO22X1 U3295 ( .IN1(n7030), .IN2(n6197), .IN3(\FIFO[36][5] ), .IN4(n6198), 
        .Q(n3384) );
  AO22X1 U3296 ( .IN1(n7019), .IN2(n6197), .IN3(\FIFO[36][6] ), .IN4(n6198), 
        .Q(n3385) );
  AO22X1 U3297 ( .IN1(n7008), .IN2(n6196), .IN3(\FIFO[36][7] ), .IN4(n6198), 
        .Q(n3386) );
  AO22X1 U3298 ( .IN1(n6997), .IN2(n6196), .IN3(\FIFO[36][8] ), .IN4(n6198), 
        .Q(n3387) );
  AO22X1 U3299 ( .IN1(n6986), .IN2(n6196), .IN3(\FIFO[36][9] ), .IN4(n6198), 
        .Q(n3388) );
  AO22X1 U3300 ( .IN1(n6975), .IN2(n6196), .IN3(\FIFO[36][10] ), .IN4(n6198), 
        .Q(n3389) );
  AO22X1 U3301 ( .IN1(n6964), .IN2(n6196), .IN3(\FIFO[36][11] ), .IN4(n6198), 
        .Q(n3390) );
  AO22X1 U3303 ( .IN1(n6942), .IN2(n6196), .IN3(\FIFO[36][13] ), .IN4(n6199), 
        .Q(n3392) );
  AO22X1 U3304 ( .IN1(n6931), .IN2(n6195), .IN3(\FIFO[36][14] ), .IN4(n6199), 
        .Q(n3393) );
  AO22X1 U3305 ( .IN1(n6920), .IN2(n6195), .IN3(\FIFO[36][15] ), .IN4(n6199), 
        .Q(n3394) );
  AO22X1 U3306 ( .IN1(n6909), .IN2(n6195), .IN3(\FIFO[36][16] ), .IN4(n6199), 
        .Q(n3395) );
  AO22X1 U3307 ( .IN1(n6898), .IN2(n6195), .IN3(\FIFO[36][17] ), .IN4(n6199), 
        .Q(n3396) );
  AO22X1 U3308 ( .IN1(n6887), .IN2(n6195), .IN3(\FIFO[36][18] ), .IN4(n6199), 
        .Q(n3397) );
  AO22X1 U3309 ( .IN1(n6876), .IN2(n6195), .IN3(\FIFO[36][19] ), .IN4(n6199), 
        .Q(n3398) );
  AO22X1 U3310 ( .IN1(n6865), .IN2(n6195), .IN3(\FIFO[36][20] ), .IN4(n6199), 
        .Q(n3399) );
  AO22X1 U3311 ( .IN1(n6854), .IN2(n6197), .IN3(\FIFO[36][21] ), .IN4(n6199), 
        .Q(n3400) );
  AO22X1 U3312 ( .IN1(n6843), .IN2(n6196), .IN3(\FIFO[36][22] ), .IN4(n6199), 
        .Q(n3401) );
  AO22X1 U3313 ( .IN1(n6832), .IN2(n6195), .IN3(\FIFO[36][23] ), .IN4(n6199), 
        .Q(n3402) );
  AO22X1 U3314 ( .IN1(n6821), .IN2(n351), .IN3(\FIFO[36][24] ), .IN4(n6200), 
        .Q(n3403) );
  AO22X1 U3315 ( .IN1(n6810), .IN2(n351), .IN3(\FIFO[36][25] ), .IN4(n6200), 
        .Q(n3404) );
  AO22X1 U3316 ( .IN1(n6799), .IN2(n351), .IN3(\FIFO[36][26] ), .IN4(n6200), 
        .Q(n3405) );
  AO22X1 U3317 ( .IN1(n6788), .IN2(n6197), .IN3(\FIFO[36][27] ), .IN4(n6200), 
        .Q(n3406) );
  AO22X1 U3318 ( .IN1(n6777), .IN2(n6196), .IN3(\FIFO[36][28] ), .IN4(n6200), 
        .Q(n3407) );
  AO22X1 U3319 ( .IN1(n6766), .IN2(n6197), .IN3(\FIFO[36][29] ), .IN4(n6200), 
        .Q(n3408) );
  AO22X1 U3320 ( .IN1(n6755), .IN2(n6196), .IN3(\FIFO[36][30] ), .IN4(n6200), 
        .Q(n3409) );
  AO22X1 U3321 ( .IN1(n6744), .IN2(n6195), .IN3(\FIFO[36][31] ), .IN4(n6200), 
        .Q(n3410) );
  AO21X1 U3322 ( .IN1(n340), .IN2(n261), .IN3(n7360), .Q(n351) );
  AO22X1 U3347 ( .IN1(n6820), .IN2(n352), .IN3(\FIFO[35][24] ), .IN4(n6194), 
        .Q(n3435) );
  AO22X1 U3348 ( .IN1(n6809), .IN2(n352), .IN3(\FIFO[35][25] ), .IN4(n6194), 
        .Q(n3436) );
  AO22X1 U3349 ( .IN1(n6798), .IN2(n352), .IN3(\FIFO[35][26] ), .IN4(n6194), 
        .Q(n3437) );
  AO22X1 U3350 ( .IN1(n6787), .IN2(n6191), .IN3(\FIFO[35][27] ), .IN4(n6194), 
        .Q(n3438) );
  AO22X1 U3351 ( .IN1(n6776), .IN2(n6191), .IN3(\FIFO[35][28] ), .IN4(n6194), 
        .Q(n3439) );
  AO22X1 U3352 ( .IN1(n6765), .IN2(n6190), .IN3(\FIFO[35][29] ), .IN4(n6194), 
        .Q(n3440) );
  AO22X1 U3353 ( .IN1(n6754), .IN2(n6189), .IN3(\FIFO[35][30] ), .IN4(n6194), 
        .Q(n3441) );
  AO22X1 U3354 ( .IN1(n6743), .IN2(n6190), .IN3(\FIFO[35][31] ), .IN4(n6194), 
        .Q(n3442) );
  AO21X1 U3355 ( .IN1(n340), .IN2(n263), .IN3(n7360), .Q(n352) );
  AO22X1 U3380 ( .IN1(n6820), .IN2(n6183), .IN3(\FIFO[34][24] ), .IN4(n6188), 
        .Q(n3467) );
  AO22X1 U3382 ( .IN1(n6798), .IN2(n6183), .IN3(\FIFO[34][26] ), .IN4(n6188), 
        .Q(n3469) );
  AO22X1 U3383 ( .IN1(n6787), .IN2(n6183), .IN3(\FIFO[34][27] ), .IN4(n6188), 
        .Q(n3470) );
  AO22X1 U3384 ( .IN1(n6776), .IN2(n6183), .IN3(\FIFO[34][28] ), .IN4(n6188), 
        .Q(n3471) );
  AO22X1 U3385 ( .IN1(n6765), .IN2(n6184), .IN3(\FIFO[34][29] ), .IN4(n6188), 
        .Q(n3472) );
  AO22X1 U3386 ( .IN1(n6754), .IN2(n6183), .IN3(\FIFO[34][30] ), .IN4(n6188), 
        .Q(n3473) );
  AO22X1 U3387 ( .IN1(n6743), .IN2(n6184), .IN3(\FIFO[34][31] ), .IN4(n6188), 
        .Q(n3474) );
  AO21X1 U3388 ( .IN1(n340), .IN2(n265), .IN3(n7360), .Q(n353) );
  AO22X1 U3389 ( .IN1(n7090), .IN2(n6179), .IN3(\FIFO[33][0] ), .IN4(n6180), 
        .Q(n3475) );
  AO22X1 U3390 ( .IN1(n7073), .IN2(n6178), .IN3(\FIFO[33][1] ), .IN4(n6180), 
        .Q(n3476) );
  AO22X1 U3391 ( .IN1(n7062), .IN2(n6177), .IN3(\FIFO[33][2] ), .IN4(n6180), 
        .Q(n3477) );
  AO22X1 U3392 ( .IN1(n7051), .IN2(n6179), .IN3(\FIFO[33][3] ), .IN4(n6180), 
        .Q(n3478) );
  AO22X1 U3393 ( .IN1(n7040), .IN2(n6178), .IN3(\FIFO[33][4] ), .IN4(n6180), 
        .Q(n3479) );
  AO22X1 U3394 ( .IN1(n7029), .IN2(n6177), .IN3(\FIFO[33][5] ), .IN4(n6180), 
        .Q(n3480) );
  AO22X1 U3395 ( .IN1(n7018), .IN2(n6179), .IN3(\FIFO[33][6] ), .IN4(n6180), 
        .Q(n3481) );
  AO22X1 U3396 ( .IN1(n7007), .IN2(n6179), .IN3(\FIFO[33][7] ), .IN4(n6180), 
        .Q(n3482) );
  AO22X1 U3397 ( .IN1(n6996), .IN2(n6179), .IN3(\FIFO[33][8] ), .IN4(n6180), 
        .Q(n3483) );
  AO22X1 U3398 ( .IN1(n6985), .IN2(n6179), .IN3(\FIFO[33][9] ), .IN4(n6180), 
        .Q(n3484) );
  AO22X1 U3399 ( .IN1(n6974), .IN2(n6179), .IN3(\FIFO[33][10] ), .IN4(n6180), 
        .Q(n3485) );
  AO22X1 U3400 ( .IN1(n6963), .IN2(n6179), .IN3(\FIFO[33][11] ), .IN4(n6180), 
        .Q(n3486) );
  AO22X1 U3401 ( .IN1(n6952), .IN2(n6179), .IN3(\FIFO[33][12] ), .IN4(n6181), 
        .Q(n3487) );
  AO22X1 U3402 ( .IN1(n6941), .IN2(n6179), .IN3(\FIFO[33][13] ), .IN4(n6181), 
        .Q(n3488) );
  AO22X1 U3403 ( .IN1(n6930), .IN2(n6178), .IN3(\FIFO[33][14] ), .IN4(n6181), 
        .Q(n3489) );
  AO22X1 U3404 ( .IN1(n6919), .IN2(n6178), .IN3(\FIFO[33][15] ), .IN4(n6181), 
        .Q(n3490) );
  AO22X1 U3405 ( .IN1(n6908), .IN2(n6178), .IN3(\FIFO[33][16] ), .IN4(n6181), 
        .Q(n3491) );
  AO22X1 U3406 ( .IN1(n6897), .IN2(n6178), .IN3(\FIFO[33][17] ), .IN4(n6181), 
        .Q(n3492) );
  AO22X1 U3408 ( .IN1(n6875), .IN2(n6178), .IN3(\FIFO[33][19] ), .IN4(n6181), 
        .Q(n3494) );
  AO22X1 U3409 ( .IN1(n6864), .IN2(n6178), .IN3(\FIFO[33][20] ), .IN4(n6181), 
        .Q(n3495) );
  AO22X1 U3410 ( .IN1(n6853), .IN2(n6177), .IN3(\FIFO[33][21] ), .IN4(n6181), 
        .Q(n3496) );
  AO22X1 U3411 ( .IN1(n6842), .IN2(n6177), .IN3(\FIFO[33][22] ), .IN4(n6181), 
        .Q(n3497) );
  AO22X1 U3412 ( .IN1(n6831), .IN2(n6177), .IN3(\FIFO[33][23] ), .IN4(n6181), 
        .Q(n3498) );
  AO22X1 U3413 ( .IN1(n6820), .IN2(n6177), .IN3(\FIFO[33][24] ), .IN4(n6182), 
        .Q(n3499) );
  AO22X1 U3414 ( .IN1(n6809), .IN2(n6177), .IN3(\FIFO[33][25] ), .IN4(n6182), 
        .Q(n3500) );
  AO22X1 U3416 ( .IN1(n6787), .IN2(n6177), .IN3(\FIFO[33][27] ), .IN4(n6182), 
        .Q(n3502) );
  AO22X1 U3417 ( .IN1(n6776), .IN2(n6177), .IN3(\FIFO[33][28] ), .IN4(n6182), 
        .Q(n3503) );
  AO22X1 U3418 ( .IN1(n6765), .IN2(n6178), .IN3(\FIFO[33][29] ), .IN4(n6182), 
        .Q(n3504) );
  AO22X1 U3419 ( .IN1(n6754), .IN2(n6177), .IN3(\FIFO[33][30] ), .IN4(n6182), 
        .Q(n3505) );
  AO22X1 U3420 ( .IN1(n6743), .IN2(n6178), .IN3(\FIFO[33][31] ), .IN4(n6182), 
        .Q(n3506) );
  AO21X1 U3421 ( .IN1(n340), .IN2(n267), .IN3(n7360), .Q(n354) );
  AO22X1 U3422 ( .IN1(n7090), .IN2(n6173), .IN3(\FIFO[32][0] ), .IN4(n6174), 
        .Q(n3507) );
  AO22X1 U3423 ( .IN1(n7073), .IN2(n6173), .IN3(\FIFO[32][1] ), .IN4(n6174), 
        .Q(n3508) );
  AO22X1 U3424 ( .IN1(n7062), .IN2(n6173), .IN3(\FIFO[32][2] ), .IN4(n6174), 
        .Q(n3509) );
  AO22X1 U3425 ( .IN1(n7051), .IN2(n6173), .IN3(\FIFO[32][3] ), .IN4(n6174), 
        .Q(n3510) );
  AO22X1 U3426 ( .IN1(n7040), .IN2(n6173), .IN3(\FIFO[32][4] ), .IN4(n6174), 
        .Q(n3511) );
  AO22X1 U3427 ( .IN1(n7029), .IN2(n6173), .IN3(\FIFO[32][5] ), .IN4(n6174), 
        .Q(n3512) );
  AO22X1 U3428 ( .IN1(n7018), .IN2(n6173), .IN3(\FIFO[32][6] ), .IN4(n6174), 
        .Q(n3513) );
  AO22X1 U3429 ( .IN1(n7007), .IN2(n6172), .IN3(\FIFO[32][7] ), .IN4(n6174), 
        .Q(n3514) );
  AO22X1 U3430 ( .IN1(n6996), .IN2(n6172), .IN3(\FIFO[32][8] ), .IN4(n6174), 
        .Q(n3515) );
  AO22X1 U3431 ( .IN1(n6985), .IN2(n6172), .IN3(\FIFO[32][9] ), .IN4(n6174), 
        .Q(n3516) );
  AO22X1 U3432 ( .IN1(n6974), .IN2(n6172), .IN3(\FIFO[32][10] ), .IN4(n6174), 
        .Q(n3517) );
  AO22X1 U3433 ( .IN1(n6963), .IN2(n6172), .IN3(\FIFO[32][11] ), .IN4(n6174), 
        .Q(n3518) );
  AO22X1 U3434 ( .IN1(n6952), .IN2(n6172), .IN3(\FIFO[32][12] ), .IN4(n6175), 
        .Q(n3519) );
  AO22X1 U3435 ( .IN1(n6941), .IN2(n6172), .IN3(\FIFO[32][13] ), .IN4(n6175), 
        .Q(n3520) );
  AO22X1 U3436 ( .IN1(n6930), .IN2(n6171), .IN3(\FIFO[32][14] ), .IN4(n6175), 
        .Q(n3521) );
  AO22X1 U3438 ( .IN1(n6908), .IN2(n6171), .IN3(\FIFO[32][16] ), .IN4(n6175), 
        .Q(n3523) );
  AO22X1 U3439 ( .IN1(n6897), .IN2(n6171), .IN3(\FIFO[32][17] ), .IN4(n6175), 
        .Q(n3524) );
  AO22X1 U3440 ( .IN1(n6886), .IN2(n6171), .IN3(\FIFO[32][18] ), .IN4(n6175), 
        .Q(n3525) );
  AO22X1 U3441 ( .IN1(n6875), .IN2(n6171), .IN3(\FIFO[32][19] ), .IN4(n6175), 
        .Q(n3526) );
  AO22X1 U3442 ( .IN1(n6864), .IN2(n6171), .IN3(\FIFO[32][20] ), .IN4(n6175), 
        .Q(n3527) );
  AO22X1 U3443 ( .IN1(n6853), .IN2(n6173), .IN3(\FIFO[32][21] ), .IN4(n6175), 
        .Q(n3528) );
  AO22X1 U3444 ( .IN1(n6842), .IN2(n6172), .IN3(\FIFO[32][22] ), .IN4(n6175), 
        .Q(n3529) );
  AO22X1 U3445 ( .IN1(n6831), .IN2(n6171), .IN3(\FIFO[32][23] ), .IN4(n6175), 
        .Q(n3530) );
  AO22X1 U3446 ( .IN1(n6820), .IN2(n355), .IN3(\FIFO[32][24] ), .IN4(n6176), 
        .Q(n3531) );
  AO22X1 U3447 ( .IN1(n6809), .IN2(n355), .IN3(\FIFO[32][25] ), .IN4(n6176), 
        .Q(n3532) );
  AO22X1 U3448 ( .IN1(n6798), .IN2(n355), .IN3(\FIFO[32][26] ), .IN4(n6176), 
        .Q(n3533) );
  AO22X1 U3449 ( .IN1(n6787), .IN2(n6173), .IN3(\FIFO[32][27] ), .IN4(n6176), 
        .Q(n3534) );
  AO22X1 U3450 ( .IN1(n6776), .IN2(n6172), .IN3(\FIFO[32][28] ), .IN4(n6176), 
        .Q(n3535) );
  AO22X1 U3451 ( .IN1(n6765), .IN2(n6173), .IN3(\FIFO[32][29] ), .IN4(n6176), 
        .Q(n3536) );
  AO22X1 U3452 ( .IN1(n6754), .IN2(n6172), .IN3(\FIFO[32][30] ), .IN4(n6176), 
        .Q(n3537) );
  AO22X1 U3453 ( .IN1(n6743), .IN2(n6171), .IN3(\FIFO[32][31] ), .IN4(n6176), 
        .Q(n3538) );
  AO21X1 U3454 ( .IN1(n340), .IN2(n269), .IN3(n7360), .Q(n355) );
  AND4X1 U3455 ( .IN1(wraddr[5]), .IN2(n270), .IN3(n7366), .IN4(n7368), .Q(
        n340) );
  AO22X1 U3480 ( .IN1(n6820), .IN2(n6165), .IN3(\FIFO[31][24] ), .IN4(n6170), 
        .Q(n3563) );
  AO22X1 U3481 ( .IN1(n6809), .IN2(n6165), .IN3(\FIFO[31][25] ), .IN4(n6170), 
        .Q(n3564) );
  AO22X1 U3482 ( .IN1(n6798), .IN2(n6165), .IN3(\FIFO[31][26] ), .IN4(n6170), 
        .Q(n3565) );
  AO22X1 U3484 ( .IN1(n6776), .IN2(n6165), .IN3(\FIFO[31][28] ), .IN4(n6170), 
        .Q(n3567) );
  AO22X1 U3485 ( .IN1(n6765), .IN2(n6166), .IN3(\FIFO[31][29] ), .IN4(n6170), 
        .Q(n3568) );
  AO22X1 U3486 ( .IN1(n6754), .IN2(n6165), .IN3(\FIFO[31][30] ), .IN4(n6170), 
        .Q(n3569) );
  AO22X1 U3487 ( .IN1(n6743), .IN2(n6166), .IN3(\FIFO[31][31] ), .IN4(n6170), 
        .Q(n3570) );
  AO21X1 U3488 ( .IN1(n357), .IN2(n238), .IN3(n7360), .Q(n356) );
  AO22X1 U3513 ( .IN1(n6820), .IN2(n358), .IN3(\FIFO[30][24] ), .IN4(n6164), 
        .Q(n3595) );
  AO22X1 U3514 ( .IN1(n6809), .IN2(n358), .IN3(\FIFO[30][25] ), .IN4(n6164), 
        .Q(n3596) );
  AO22X1 U3515 ( .IN1(n6798), .IN2(n358), .IN3(\FIFO[30][26] ), .IN4(n6164), 
        .Q(n3597) );
  AO22X1 U3516 ( .IN1(n6787), .IN2(n6161), .IN3(\FIFO[30][27] ), .IN4(n6164), 
        .Q(n3598) );
  AO22X1 U3517 ( .IN1(n6776), .IN2(n6160), .IN3(\FIFO[30][28] ), .IN4(n6164), 
        .Q(n3599) );
  AO22X1 U3518 ( .IN1(n6765), .IN2(n6161), .IN3(\FIFO[30][29] ), .IN4(n6164), 
        .Q(n3600) );
  AO22X1 U3519 ( .IN1(n6754), .IN2(n6160), .IN3(\FIFO[30][30] ), .IN4(n6164), 
        .Q(n3601) );
  AO22X1 U3520 ( .IN1(n6743), .IN2(n6159), .IN3(\FIFO[30][31] ), .IN4(n6164), 
        .Q(n3602) );
  AO21X1 U3521 ( .IN1(n357), .IN2(n241), .IN3(n7360), .Q(n358) );
  AO22X1 U3522 ( .IN1(n7090), .IN2(n6155), .IN3(\FIFO[29][0] ), .IN4(n6156), 
        .Q(n3603) );
  AO22X1 U3523 ( .IN1(n7073), .IN2(n6155), .IN3(\FIFO[29][1] ), .IN4(n6156), 
        .Q(n3604) );
  AO22X1 U3525 ( .IN1(n7051), .IN2(n6155), .IN3(\FIFO[29][3] ), .IN4(n6156), 
        .Q(n3606) );
  AO22X1 U3526 ( .IN1(n7040), .IN2(n6155), .IN3(\FIFO[29][4] ), .IN4(n6156), 
        .Q(n3607) );
  AO22X1 U3527 ( .IN1(n7029), .IN2(n6155), .IN3(\FIFO[29][5] ), .IN4(n6156), 
        .Q(n3608) );
  AO22X1 U3528 ( .IN1(n7018), .IN2(n6155), .IN3(\FIFO[29][6] ), .IN4(n6156), 
        .Q(n3609) );
  AO22X1 U3529 ( .IN1(n7007), .IN2(n6154), .IN3(\FIFO[29][7] ), .IN4(n6156), 
        .Q(n3610) );
  AO22X1 U3530 ( .IN1(n6996), .IN2(n6154), .IN3(\FIFO[29][8] ), .IN4(n6156), 
        .Q(n3611) );
  AO22X1 U3531 ( .IN1(n6985), .IN2(n6154), .IN3(\FIFO[29][9] ), .IN4(n6156), 
        .Q(n3612) );
  AO22X1 U3532 ( .IN1(n6974), .IN2(n6154), .IN3(\FIFO[29][10] ), .IN4(n6156), 
        .Q(n3613) );
  AO22X1 U3533 ( .IN1(n6963), .IN2(n6154), .IN3(\FIFO[29][11] ), .IN4(n6156), 
        .Q(n3614) );
  AO22X1 U3534 ( .IN1(n6952), .IN2(n6154), .IN3(\FIFO[29][12] ), .IN4(n6157), 
        .Q(n3615) );
  AO22X1 U3535 ( .IN1(n6941), .IN2(n6154), .IN3(\FIFO[29][13] ), .IN4(n6157), 
        .Q(n3616) );
  AO22X1 U3536 ( .IN1(n6930), .IN2(n6153), .IN3(\FIFO[29][14] ), .IN4(n6157), 
        .Q(n3617) );
  AO22X1 U3537 ( .IN1(n6919), .IN2(n6153), .IN3(\FIFO[29][15] ), .IN4(n6157), 
        .Q(n3618) );
  AO22X1 U3538 ( .IN1(n6908), .IN2(n6153), .IN3(\FIFO[29][16] ), .IN4(n6157), 
        .Q(n3619) );
  AO22X1 U3539 ( .IN1(n6897), .IN2(n6153), .IN3(\FIFO[29][17] ), .IN4(n6157), 
        .Q(n3620) );
  AO22X1 U3540 ( .IN1(n6886), .IN2(n6153), .IN3(\FIFO[29][18] ), .IN4(n6157), 
        .Q(n3621) );
  AO22X1 U3541 ( .IN1(n6875), .IN2(n6153), .IN3(\FIFO[29][19] ), .IN4(n6157), 
        .Q(n3622) );
  AO22X1 U3542 ( .IN1(n6864), .IN2(n6153), .IN3(\FIFO[29][20] ), .IN4(n6157), 
        .Q(n3623) );
  AO22X1 U3543 ( .IN1(n6853), .IN2(n6155), .IN3(\FIFO[29][21] ), .IN4(n6157), 
        .Q(n3624) );
  AO22X1 U3544 ( .IN1(n6842), .IN2(n6154), .IN3(\FIFO[29][22] ), .IN4(n6157), 
        .Q(n3625) );
  AO22X1 U3545 ( .IN1(n6831), .IN2(n6153), .IN3(\FIFO[29][23] ), .IN4(n6157), 
        .Q(n3626) );
  AO22X1 U3546 ( .IN1(n6820), .IN2(n359), .IN3(\FIFO[29][24] ), .IN4(n6158), 
        .Q(n3627) );
  AO22X1 U3547 ( .IN1(n6809), .IN2(n359), .IN3(\FIFO[29][25] ), .IN4(n6158), 
        .Q(n3628) );
  AO22X1 U3548 ( .IN1(n6798), .IN2(n359), .IN3(\FIFO[29][26] ), .IN4(n6158), 
        .Q(n3629) );
  AO22X1 U3549 ( .IN1(n6787), .IN2(n6155), .IN3(\FIFO[29][27] ), .IN4(n6158), 
        .Q(n3630) );
  AO22X1 U3550 ( .IN1(n6776), .IN2(n6154), .IN3(\FIFO[29][28] ), .IN4(n6158), 
        .Q(n3631) );
  AO22X1 U3551 ( .IN1(n6765), .IN2(n6155), .IN3(\FIFO[29][29] ), .IN4(n6158), 
        .Q(n3632) );
  AO22X1 U3552 ( .IN1(n6754), .IN2(n6154), .IN3(\FIFO[29][30] ), .IN4(n6158), 
        .Q(n3633) );
  AO22X1 U3553 ( .IN1(n6743), .IN2(n6153), .IN3(\FIFO[29][31] ), .IN4(n6158), 
        .Q(n3634) );
  AO21X1 U3554 ( .IN1(n357), .IN2(n243), .IN3(n7360), .Q(n359) );
  AO22X1 U3555 ( .IN1(n7090), .IN2(n6149), .IN3(\FIFO[28][0] ), .IN4(n6150), 
        .Q(n3635) );
  AO22X1 U3556 ( .IN1(n7073), .IN2(n6149), .IN3(\FIFO[28][1] ), .IN4(n6150), 
        .Q(n3636) );
  AO22X1 U3557 ( .IN1(n7062), .IN2(n6149), .IN3(\FIFO[28][2] ), .IN4(n6150), 
        .Q(n3637) );
  AO22X1 U3559 ( .IN1(n7040), .IN2(n6149), .IN3(\FIFO[28][4] ), .IN4(n6150), 
        .Q(n3639) );
  AO22X1 U3560 ( .IN1(n7029), .IN2(n6149), .IN3(\FIFO[28][5] ), .IN4(n6150), 
        .Q(n3640) );
  AO22X1 U3561 ( .IN1(n7018), .IN2(n6149), .IN3(\FIFO[28][6] ), .IN4(n6150), 
        .Q(n3641) );
  AO22X1 U3562 ( .IN1(n7007), .IN2(n6148), .IN3(\FIFO[28][7] ), .IN4(n6150), 
        .Q(n3642) );
  AO22X1 U3563 ( .IN1(n6996), .IN2(n6148), .IN3(\FIFO[28][8] ), .IN4(n6150), 
        .Q(n3643) );
  AO22X1 U3564 ( .IN1(n6985), .IN2(n6148), .IN3(\FIFO[28][9] ), .IN4(n6150), 
        .Q(n3644) );
  AO22X1 U3565 ( .IN1(n6974), .IN2(n6148), .IN3(\FIFO[28][10] ), .IN4(n6150), 
        .Q(n3645) );
  AO22X1 U3566 ( .IN1(n6963), .IN2(n6148), .IN3(\FIFO[28][11] ), .IN4(n6150), 
        .Q(n3646) );
  AO22X1 U3568 ( .IN1(n6941), .IN2(n6148), .IN3(\FIFO[28][13] ), .IN4(n6151), 
        .Q(n3648) );
  AO22X1 U3569 ( .IN1(n6930), .IN2(n6147), .IN3(\FIFO[28][14] ), .IN4(n6151), 
        .Q(n3649) );
  AO22X1 U3570 ( .IN1(n6919), .IN2(n6147), .IN3(\FIFO[28][15] ), .IN4(n6151), 
        .Q(n3650) );
  AO22X1 U3571 ( .IN1(n6908), .IN2(n6147), .IN3(\FIFO[28][16] ), .IN4(n6151), 
        .Q(n3651) );
  AO22X1 U3572 ( .IN1(n6897), .IN2(n6147), .IN3(\FIFO[28][17] ), .IN4(n6151), 
        .Q(n3652) );
  AO22X1 U3573 ( .IN1(n6886), .IN2(n6147), .IN3(\FIFO[28][18] ), .IN4(n6151), 
        .Q(n3653) );
  AO22X1 U3574 ( .IN1(n6875), .IN2(n6147), .IN3(\FIFO[28][19] ), .IN4(n6151), 
        .Q(n3654) );
  AO22X1 U3575 ( .IN1(n6864), .IN2(n6147), .IN3(\FIFO[28][20] ), .IN4(n6151), 
        .Q(n3655) );
  AO22X1 U3576 ( .IN1(n6853), .IN2(n6149), .IN3(\FIFO[28][21] ), .IN4(n6151), 
        .Q(n3656) );
  AO22X1 U3577 ( .IN1(n6842), .IN2(n6148), .IN3(\FIFO[28][22] ), .IN4(n6151), 
        .Q(n3657) );
  AO22X1 U3578 ( .IN1(n6831), .IN2(n6147), .IN3(\FIFO[28][23] ), .IN4(n6151), 
        .Q(n3658) );
  AO22X1 U3579 ( .IN1(n6820), .IN2(n360), .IN3(\FIFO[28][24] ), .IN4(n6152), 
        .Q(n3659) );
  AO22X1 U3580 ( .IN1(n6809), .IN2(n360), .IN3(\FIFO[28][25] ), .IN4(n6152), 
        .Q(n3660) );
  AO22X1 U3581 ( .IN1(n6798), .IN2(n360), .IN3(\FIFO[28][26] ), .IN4(n6152), 
        .Q(n3661) );
  AO22X1 U3582 ( .IN1(n6787), .IN2(n6149), .IN3(\FIFO[28][27] ), .IN4(n6152), 
        .Q(n3662) );
  AO22X1 U3583 ( .IN1(n6776), .IN2(n6149), .IN3(\FIFO[28][28] ), .IN4(n6152), 
        .Q(n3663) );
  AO22X1 U3584 ( .IN1(n6765), .IN2(n6148), .IN3(\FIFO[28][29] ), .IN4(n6152), 
        .Q(n3664) );
  AO22X1 U3585 ( .IN1(n6754), .IN2(n6147), .IN3(\FIFO[28][30] ), .IN4(n6152), 
        .Q(n3665) );
  AO22X1 U3586 ( .IN1(n6743), .IN2(n6148), .IN3(\FIFO[28][31] ), .IN4(n6152), 
        .Q(n3666) );
  AO21X1 U3587 ( .IN1(n357), .IN2(n245), .IN3(n7360), .Q(n360) );
  AO22X1 U3612 ( .IN1(n6820), .IN2(n6141), .IN3(\FIFO[27][24] ), .IN4(n6146), 
        .Q(n3691) );
  AO22X1 U3613 ( .IN1(n6809), .IN2(n6141), .IN3(\FIFO[27][25] ), .IN4(n6146), 
        .Q(n3692) );
  AO22X1 U3614 ( .IN1(n6798), .IN2(n6141), .IN3(\FIFO[27][26] ), .IN4(n6146), 
        .Q(n3693) );
  AO22X1 U3615 ( .IN1(n6787), .IN2(n6141), .IN3(\FIFO[27][27] ), .IN4(n6146), 
        .Q(n3694) );
  AO22X1 U3617 ( .IN1(n6765), .IN2(n6142), .IN3(\FIFO[27][29] ), .IN4(n6146), 
        .Q(n3696) );
  AO22X1 U3618 ( .IN1(n6754), .IN2(n6141), .IN3(\FIFO[27][30] ), .IN4(n6146), 
        .Q(n3697) );
  AO22X1 U3619 ( .IN1(n6743), .IN2(n6142), .IN3(\FIFO[27][31] ), .IN4(n6146), 
        .Q(n3698) );
  AO21X1 U3620 ( .IN1(n357), .IN2(n247), .IN3(n7360), .Q(n361) );
  AO22X1 U3645 ( .IN1(n6820), .IN2(n6135), .IN3(\FIFO[26][24] ), .IN4(n6140), 
        .Q(n3723) );
  AO22X1 U3646 ( .IN1(n6809), .IN2(n6135), .IN3(\FIFO[26][25] ), .IN4(n6140), 
        .Q(n3724) );
  AO22X1 U3647 ( .IN1(n6798), .IN2(n6135), .IN3(\FIFO[26][26] ), .IN4(n6140), 
        .Q(n3725) );
  AO22X1 U3648 ( .IN1(n6787), .IN2(n6135), .IN3(\FIFO[26][27] ), .IN4(n6140), 
        .Q(n3726) );
  AO22X1 U3649 ( .IN1(n6776), .IN2(n6135), .IN3(\FIFO[26][28] ), .IN4(n6140), 
        .Q(n3727) );
  AO22X1 U3651 ( .IN1(n6754), .IN2(n6135), .IN3(\FIFO[26][30] ), .IN4(n6140), 
        .Q(n3729) );
  AO22X1 U3652 ( .IN1(n6743), .IN2(n6136), .IN3(\FIFO[26][31] ), .IN4(n6140), 
        .Q(n3730) );
  AO21X1 U3653 ( .IN1(n357), .IN2(n249), .IN3(n7360), .Q(n362) );
  AO22X1 U3654 ( .IN1(n7090), .IN2(n6131), .IN3(\FIFO[25][0] ), .IN4(n6132), 
        .Q(n3731) );
  AO22X1 U3655 ( .IN1(n7073), .IN2(n6131), .IN3(\FIFO[25][1] ), .IN4(n6132), 
        .Q(n3732) );
  AO22X1 U3656 ( .IN1(n7062), .IN2(n6131), .IN3(\FIFO[25][2] ), .IN4(n6132), 
        .Q(n3733) );
  AO22X1 U3657 ( .IN1(n7051), .IN2(n6131), .IN3(\FIFO[25][3] ), .IN4(n6132), 
        .Q(n3734) );
  AO22X1 U3658 ( .IN1(n7040), .IN2(n6131), .IN3(\FIFO[25][4] ), .IN4(n6132), 
        .Q(n3735) );
  AO22X1 U3659 ( .IN1(n7029), .IN2(n6131), .IN3(\FIFO[25][5] ), .IN4(n6132), 
        .Q(n3736) );
  AO22X1 U3661 ( .IN1(n7007), .IN2(n6130), .IN3(\FIFO[25][7] ), .IN4(n6132), 
        .Q(n3738) );
  AO22X1 U3662 ( .IN1(n6996), .IN2(n6130), .IN3(\FIFO[25][8] ), .IN4(n6132), 
        .Q(n3739) );
  AO22X1 U3663 ( .IN1(n6985), .IN2(n6130), .IN3(\FIFO[25][9] ), .IN4(n6132), 
        .Q(n3740) );
  AO22X1 U3664 ( .IN1(n6974), .IN2(n6130), .IN3(\FIFO[25][10] ), .IN4(n6132), 
        .Q(n3741) );
  AO22X1 U3665 ( .IN1(n6963), .IN2(n6130), .IN3(\FIFO[25][11] ), .IN4(n6132), 
        .Q(n3742) );
  AO22X1 U3666 ( .IN1(n6952), .IN2(n6130), .IN3(\FIFO[25][12] ), .IN4(n6133), 
        .Q(n3743) );
  AO22X1 U3668 ( .IN1(n6930), .IN2(n6129), .IN3(\FIFO[25][14] ), .IN4(n6133), 
        .Q(n3745) );
  AO22X1 U3669 ( .IN1(n6919), .IN2(n6129), .IN3(\FIFO[25][15] ), .IN4(n6133), 
        .Q(n3746) );
  AO22X1 U3670 ( .IN1(n6908), .IN2(n6129), .IN3(\FIFO[25][16] ), .IN4(n6133), 
        .Q(n3747) );
  AO22X1 U3671 ( .IN1(n6897), .IN2(n6129), .IN3(\FIFO[25][17] ), .IN4(n6133), 
        .Q(n3748) );
  AO22X1 U3672 ( .IN1(n6886), .IN2(n6129), .IN3(\FIFO[25][18] ), .IN4(n6133), 
        .Q(n3749) );
  AO22X1 U3673 ( .IN1(n6875), .IN2(n6129), .IN3(\FIFO[25][19] ), .IN4(n6133), 
        .Q(n3750) );
  AO22X1 U3674 ( .IN1(n6864), .IN2(n6129), .IN3(\FIFO[25][20] ), .IN4(n6133), 
        .Q(n3751) );
  AO22X1 U3675 ( .IN1(n6853), .IN2(n6131), .IN3(\FIFO[25][21] ), .IN4(n6133), 
        .Q(n3752) );
  AO22X1 U3676 ( .IN1(n6842), .IN2(n6130), .IN3(\FIFO[25][22] ), .IN4(n6133), 
        .Q(n3753) );
  AO22X1 U3677 ( .IN1(n6831), .IN2(n6129), .IN3(\FIFO[25][23] ), .IN4(n6133), 
        .Q(n3754) );
  AO22X1 U3678 ( .IN1(n6820), .IN2(n363), .IN3(\FIFO[25][24] ), .IN4(n6134), 
        .Q(n3755) );
  AO22X1 U3679 ( .IN1(n6809), .IN2(n363), .IN3(\FIFO[25][25] ), .IN4(n6134), 
        .Q(n3756) );
  AO22X1 U3680 ( .IN1(n6798), .IN2(n363), .IN3(\FIFO[25][26] ), .IN4(n6134), 
        .Q(n3757) );
  AO22X1 U3681 ( .IN1(n6787), .IN2(n6131), .IN3(\FIFO[25][27] ), .IN4(n6134), 
        .Q(n3758) );
  AO22X1 U3682 ( .IN1(n6776), .IN2(n6130), .IN3(\FIFO[25][28] ), .IN4(n6134), 
        .Q(n3759) );
  AO22X1 U3683 ( .IN1(n6765), .IN2(n6131), .IN3(\FIFO[25][29] ), .IN4(n6134), 
        .Q(n3760) );
  AO22X1 U3684 ( .IN1(n6754), .IN2(n6130), .IN3(\FIFO[25][30] ), .IN4(n6134), 
        .Q(n3761) );
  AO22X1 U3685 ( .IN1(n6743), .IN2(n6129), .IN3(\FIFO[25][31] ), .IN4(n6134), 
        .Q(n3762) );
  AO21X1 U3686 ( .IN1(n357), .IN2(n251), .IN3(n7361), .Q(n363) );
  AO22X1 U3687 ( .IN1(n7090), .IN2(n6125), .IN3(\FIFO[24][0] ), .IN4(n6126), 
        .Q(n3763) );
  AO22X1 U3688 ( .IN1(n7073), .IN2(n6125), .IN3(\FIFO[24][1] ), .IN4(n6126), 
        .Q(n3764) );
  AO22X1 U3689 ( .IN1(n7062), .IN2(n6125), .IN3(\FIFO[24][2] ), .IN4(n6126), 
        .Q(n3765) );
  AO22X1 U3690 ( .IN1(n7051), .IN2(n6125), .IN3(\FIFO[24][3] ), .IN4(n6126), 
        .Q(n3766) );
  AO22X1 U3691 ( .IN1(n7040), .IN2(n6125), .IN3(\FIFO[24][4] ), .IN4(n6126), 
        .Q(n3767) );
  AO22X1 U3692 ( .IN1(n7029), .IN2(n6125), .IN3(\FIFO[24][5] ), .IN4(n6126), 
        .Q(n3768) );
  AO22X1 U3693 ( .IN1(n7018), .IN2(n6125), .IN3(\FIFO[24][6] ), .IN4(n6126), 
        .Q(n3769) );
  AO22X1 U3695 ( .IN1(n6996), .IN2(n6124), .IN3(\FIFO[24][8] ), .IN4(n6126), 
        .Q(n3771) );
  AO22X1 U3696 ( .IN1(n6985), .IN2(n6124), .IN3(\FIFO[24][9] ), .IN4(n6126), 
        .Q(n3772) );
  AO22X1 U3697 ( .IN1(n6974), .IN2(n6124), .IN3(\FIFO[24][10] ), .IN4(n6126), 
        .Q(n3773) );
  AO22X1 U3698 ( .IN1(n6963), .IN2(n6124), .IN3(\FIFO[24][11] ), .IN4(n6126), 
        .Q(n3774) );
  AO22X1 U3699 ( .IN1(n6952), .IN2(n6124), .IN3(\FIFO[24][12] ), .IN4(n6127), 
        .Q(n3775) );
  AO22X1 U3700 ( .IN1(n6941), .IN2(n6124), .IN3(\FIFO[24][13] ), .IN4(n6127), 
        .Q(n3776) );
  AO22X1 U3701 ( .IN1(n6930), .IN2(n6123), .IN3(\FIFO[24][14] ), .IN4(n6127), 
        .Q(n3777) );
  AO22X1 U3702 ( .IN1(n6919), .IN2(n6123), .IN3(\FIFO[24][15] ), .IN4(n6127), 
        .Q(n3778) );
  AO22X1 U3703 ( .IN1(n6908), .IN2(n6123), .IN3(\FIFO[24][16] ), .IN4(n6127), 
        .Q(n3779) );
  AO22X1 U3704 ( .IN1(n6897), .IN2(n6123), .IN3(\FIFO[24][17] ), .IN4(n6127), 
        .Q(n3780) );
  AO22X1 U3705 ( .IN1(n6886), .IN2(n6123), .IN3(\FIFO[24][18] ), .IN4(n6127), 
        .Q(n3781) );
  AO22X1 U3706 ( .IN1(n6875), .IN2(n6123), .IN3(\FIFO[24][19] ), .IN4(n6127), 
        .Q(n3782) );
  AO22X1 U3707 ( .IN1(n6864), .IN2(n6123), .IN3(\FIFO[24][20] ), .IN4(n6127), 
        .Q(n3783) );
  AO22X1 U3708 ( .IN1(n6853), .IN2(n6125), .IN3(\FIFO[24][21] ), .IN4(n6127), 
        .Q(n3784) );
  AO22X1 U3709 ( .IN1(n6842), .IN2(n6124), .IN3(\FIFO[24][22] ), .IN4(n6127), 
        .Q(n3785) );
  AO22X1 U3710 ( .IN1(n6831), .IN2(n6123), .IN3(\FIFO[24][23] ), .IN4(n6127), 
        .Q(n3786) );
  AO22X1 U3711 ( .IN1(n6820), .IN2(n364), .IN3(\FIFO[24][24] ), .IN4(n6128), 
        .Q(n3787) );
  AO22X1 U3712 ( .IN1(n6809), .IN2(n364), .IN3(\FIFO[24][25] ), .IN4(n6128), 
        .Q(n3788) );
  AO22X1 U3713 ( .IN1(n6798), .IN2(n364), .IN3(\FIFO[24][26] ), .IN4(n6128), 
        .Q(n3789) );
  AO22X1 U3714 ( .IN1(n6787), .IN2(n6125), .IN3(\FIFO[24][27] ), .IN4(n6128), 
        .Q(n3790) );
  AO22X1 U3715 ( .IN1(n6776), .IN2(n6124), .IN3(\FIFO[24][28] ), .IN4(n6128), 
        .Q(n3791) );
  AO22X1 U3716 ( .IN1(n6765), .IN2(n6125), .IN3(\FIFO[24][29] ), .IN4(n6128), 
        .Q(n3792) );
  AO22X1 U3717 ( .IN1(n6754), .IN2(n6124), .IN3(\FIFO[24][30] ), .IN4(n6128), 
        .Q(n3793) );
  AO22X1 U3718 ( .IN1(n6743), .IN2(n6123), .IN3(\FIFO[24][31] ), .IN4(n6128), 
        .Q(n3794) );
  AO21X1 U3719 ( .IN1(n357), .IN2(n253), .IN3(n7361), .Q(n364) );
  AO22X1 U3744 ( .IN1(n6819), .IN2(n365), .IN3(\FIFO[23][24] ), .IN4(n6122), 
        .Q(n3819) );
  AO22X1 U3745 ( .IN1(n6808), .IN2(n365), .IN3(\FIFO[23][25] ), .IN4(n6122), 
        .Q(n3820) );
  AO22X1 U3746 ( .IN1(n6797), .IN2(n365), .IN3(\FIFO[23][26] ), .IN4(n6122), 
        .Q(n3821) );
  AO22X1 U3747 ( .IN1(n6786), .IN2(n6119), .IN3(\FIFO[23][27] ), .IN4(n6122), 
        .Q(n3822) );
  AO22X1 U3748 ( .IN1(n6775), .IN2(n6119), .IN3(\FIFO[23][28] ), .IN4(n6122), 
        .Q(n3823) );
  AO22X1 U3749 ( .IN1(n6764), .IN2(n6118), .IN3(\FIFO[23][29] ), .IN4(n6122), 
        .Q(n3824) );
  AO22X1 U3750 ( .IN1(n6753), .IN2(n6117), .IN3(\FIFO[23][30] ), .IN4(n6122), 
        .Q(n3825) );
  AO22X1 U3751 ( .IN1(n6742), .IN2(n6118), .IN3(\FIFO[23][31] ), .IN4(n6122), 
        .Q(n3826) );
  AO21X1 U3752 ( .IN1(n357), .IN2(n255), .IN3(n7361), .Q(n365) );
  AO22X1 U3777 ( .IN1(n6819), .IN2(n6111), .IN3(\FIFO[22][24] ), .IN4(n6116), 
        .Q(n3851) );
  AO22X1 U3778 ( .IN1(n6808), .IN2(n6111), .IN3(\FIFO[22][25] ), .IN4(n6116), 
        .Q(n3852) );
  AO22X1 U3779 ( .IN1(n6797), .IN2(n6111), .IN3(\FIFO[22][26] ), .IN4(n6116), 
        .Q(n3853) );
  AO22X1 U3780 ( .IN1(n6786), .IN2(n6111), .IN3(\FIFO[22][27] ), .IN4(n6116), 
        .Q(n3854) );
  AO22X1 U3781 ( .IN1(n6775), .IN2(n6111), .IN3(\FIFO[22][28] ), .IN4(n6116), 
        .Q(n3855) );
  AO22X1 U3782 ( .IN1(n6764), .IN2(n6112), .IN3(\FIFO[22][29] ), .IN4(n6116), 
        .Q(n3856) );
  AO22X1 U3784 ( .IN1(n6742), .IN2(n6112), .IN3(\FIFO[22][31] ), .IN4(n6116), 
        .Q(n3858) );
  AO21X1 U3785 ( .IN1(n357), .IN2(n257), .IN3(n7361), .Q(n366) );
  AO22X1 U3786 ( .IN1(n7089), .IN2(n6107), .IN3(\FIFO[21][0] ), .IN4(n6108), 
        .Q(n3859) );
  AO22X1 U3787 ( .IN1(n7072), .IN2(n6106), .IN3(\FIFO[21][1] ), .IN4(n6108), 
        .Q(n3860) );
  AO22X1 U3788 ( .IN1(n7061), .IN2(n6105), .IN3(\FIFO[21][2] ), .IN4(n6108), 
        .Q(n3861) );
  AO22X1 U3789 ( .IN1(n7050), .IN2(n6107), .IN3(\FIFO[21][3] ), .IN4(n6108), 
        .Q(n3862) );
  AO22X1 U3790 ( .IN1(n7039), .IN2(n6106), .IN3(\FIFO[21][4] ), .IN4(n6108), 
        .Q(n3863) );
  AO22X1 U3791 ( .IN1(n7028), .IN2(n6105), .IN3(\FIFO[21][5] ), .IN4(n6108), 
        .Q(n3864) );
  AO22X1 U3792 ( .IN1(n7017), .IN2(n6107), .IN3(\FIFO[21][6] ), .IN4(n6108), 
        .Q(n3865) );
  AO22X1 U3793 ( .IN1(n7006), .IN2(n6107), .IN3(\FIFO[21][7] ), .IN4(n6108), 
        .Q(n3866) );
  AO22X1 U3794 ( .IN1(n6995), .IN2(n6107), .IN3(\FIFO[21][8] ), .IN4(n6108), 
        .Q(n3867) );
  AO22X1 U3795 ( .IN1(n6984), .IN2(n6107), .IN3(\FIFO[21][9] ), .IN4(n6108), 
        .Q(n3868) );
  AO22X1 U3797 ( .IN1(n6962), .IN2(n6107), .IN3(\FIFO[21][11] ), .IN4(n6108), 
        .Q(n3870) );
  AO22X1 U3798 ( .IN1(n6951), .IN2(n6107), .IN3(\FIFO[21][12] ), .IN4(n6109), 
        .Q(n3871) );
  AO22X1 U3799 ( .IN1(n6940), .IN2(n6107), .IN3(\FIFO[21][13] ), .IN4(n6109), 
        .Q(n3872) );
  AO22X1 U3800 ( .IN1(n6929), .IN2(n6106), .IN3(\FIFO[21][14] ), .IN4(n6109), 
        .Q(n3873) );
  AO22X1 U3801 ( .IN1(n6918), .IN2(n6106), .IN3(\FIFO[21][15] ), .IN4(n6109), 
        .Q(n3874) );
  AO22X1 U3802 ( .IN1(n6907), .IN2(n6106), .IN3(\FIFO[21][16] ), .IN4(n6109), 
        .Q(n3875) );
  AO22X1 U3803 ( .IN1(n6896), .IN2(n6106), .IN3(\FIFO[21][17] ), .IN4(n6109), 
        .Q(n3876) );
  AO22X1 U3804 ( .IN1(n6885), .IN2(n6106), .IN3(\FIFO[21][18] ), .IN4(n6109), 
        .Q(n3877) );
  AO22X1 U3805 ( .IN1(n6874), .IN2(n6106), .IN3(\FIFO[21][19] ), .IN4(n6109), 
        .Q(n3878) );
  AO22X1 U3806 ( .IN1(n6863), .IN2(n6106), .IN3(\FIFO[21][20] ), .IN4(n6109), 
        .Q(n3879) );
  AO22X1 U3807 ( .IN1(n6852), .IN2(n6105), .IN3(\FIFO[21][21] ), .IN4(n6109), 
        .Q(n3880) );
  AO22X1 U3808 ( .IN1(n6841), .IN2(n6105), .IN3(\FIFO[21][22] ), .IN4(n6109), 
        .Q(n3881) );
  AO22X1 U3810 ( .IN1(n6819), .IN2(n6105), .IN3(\FIFO[21][24] ), .IN4(n6110), 
        .Q(n3883) );
  AO22X1 U3811 ( .IN1(n6808), .IN2(n6105), .IN3(\FIFO[21][25] ), .IN4(n6110), 
        .Q(n3884) );
  AO22X1 U3812 ( .IN1(n6797), .IN2(n6105), .IN3(\FIFO[21][26] ), .IN4(n6110), 
        .Q(n3885) );
  AO22X1 U3813 ( .IN1(n6786), .IN2(n6105), .IN3(\FIFO[21][27] ), .IN4(n6110), 
        .Q(n3886) );
  AO22X1 U3814 ( .IN1(n6775), .IN2(n6105), .IN3(\FIFO[21][28] ), .IN4(n6110), 
        .Q(n3887) );
  AO22X1 U3815 ( .IN1(n6764), .IN2(n6106), .IN3(\FIFO[21][29] ), .IN4(n6110), 
        .Q(n3888) );
  AO22X1 U3816 ( .IN1(n6753), .IN2(n6105), .IN3(\FIFO[21][30] ), .IN4(n6110), 
        .Q(n3889) );
  AO21X1 U3818 ( .IN1(n357), .IN2(n259), .IN3(n7361), .Q(n367) );
  AO22X1 U3819 ( .IN1(n7089), .IN2(n6101), .IN3(\FIFO[20][0] ), .IN4(n6102), 
        .Q(n3891) );
  AO22X1 U3820 ( .IN1(n7072), .IN2(n6101), .IN3(\FIFO[20][1] ), .IN4(n6102), 
        .Q(n3892) );
  AO22X1 U3821 ( .IN1(n7061), .IN2(n6101), .IN3(\FIFO[20][2] ), .IN4(n6102), 
        .Q(n3893) );
  AO22X1 U3822 ( .IN1(n7050), .IN2(n6101), .IN3(\FIFO[20][3] ), .IN4(n6102), 
        .Q(n3894) );
  AO22X1 U3823 ( .IN1(n7039), .IN2(n6101), .IN3(\FIFO[20][4] ), .IN4(n6102), 
        .Q(n3895) );
  AO22X1 U3824 ( .IN1(n7028), .IN2(n6101), .IN3(\FIFO[20][5] ), .IN4(n6102), 
        .Q(n3896) );
  AO22X1 U3825 ( .IN1(n7017), .IN2(n6101), .IN3(\FIFO[20][6] ), .IN4(n6102), 
        .Q(n3897) );
  AO22X1 U3826 ( .IN1(n7006), .IN2(n6100), .IN3(\FIFO[20][7] ), .IN4(n6102), 
        .Q(n3898) );
  AO22X1 U3827 ( .IN1(n6995), .IN2(n6100), .IN3(\FIFO[20][8] ), .IN4(n6102), 
        .Q(n3899) );
  AO22X1 U3828 ( .IN1(n6984), .IN2(n6100), .IN3(\FIFO[20][9] ), .IN4(n6102), 
        .Q(n3900) );
  AO22X1 U3829 ( .IN1(n6973), .IN2(n6100), .IN3(\FIFO[20][10] ), .IN4(n6102), 
        .Q(n3901) );
  AO22X1 U3831 ( .IN1(n6951), .IN2(n6100), .IN3(\FIFO[20][12] ), .IN4(n6103), 
        .Q(n3903) );
  AO22X1 U3832 ( .IN1(n6940), .IN2(n6100), .IN3(\FIFO[20][13] ), .IN4(n6103), 
        .Q(n3904) );
  AO22X1 U3833 ( .IN1(n6929), .IN2(n6099), .IN3(\FIFO[20][14] ), .IN4(n6103), 
        .Q(n3905) );
  AO22X1 U3834 ( .IN1(n6918), .IN2(n6099), .IN3(\FIFO[20][15] ), .IN4(n6103), 
        .Q(n3906) );
  AO22X1 U3835 ( .IN1(n6907), .IN2(n6099), .IN3(\FIFO[20][16] ), .IN4(n6103), 
        .Q(n3907) );
  AO22X1 U3836 ( .IN1(n6896), .IN2(n6099), .IN3(\FIFO[20][17] ), .IN4(n6103), 
        .Q(n3908) );
  AO22X1 U3837 ( .IN1(n6885), .IN2(n6099), .IN3(\FIFO[20][18] ), .IN4(n6103), 
        .Q(n3909) );
  AO22X1 U3838 ( .IN1(n6874), .IN2(n6099), .IN3(\FIFO[20][19] ), .IN4(n6103), 
        .Q(n3910) );
  AO22X1 U3839 ( .IN1(n6863), .IN2(n6099), .IN3(\FIFO[20][20] ), .IN4(n6103), 
        .Q(n3911) );
  AO22X1 U3840 ( .IN1(n6852), .IN2(n6101), .IN3(\FIFO[20][21] ), .IN4(n6103), 
        .Q(n3912) );
  AO22X1 U3841 ( .IN1(n6841), .IN2(n6100), .IN3(\FIFO[20][22] ), .IN4(n6103), 
        .Q(n3913) );
  AO22X1 U3842 ( .IN1(n6830), .IN2(n6099), .IN3(\FIFO[20][23] ), .IN4(n6103), 
        .Q(n3914) );
  AO22X1 U3843 ( .IN1(n6819), .IN2(n368), .IN3(\FIFO[20][24] ), .IN4(n6104), 
        .Q(n3915) );
  AO22X1 U3844 ( .IN1(n6808), .IN2(n368), .IN3(\FIFO[20][25] ), .IN4(n6104), 
        .Q(n3916) );
  AO22X1 U3845 ( .IN1(n6797), .IN2(n368), .IN3(\FIFO[20][26] ), .IN4(n6104), 
        .Q(n3917) );
  AO22X1 U3846 ( .IN1(n6786), .IN2(n6101), .IN3(\FIFO[20][27] ), .IN4(n6104), 
        .Q(n3918) );
  AO22X1 U3847 ( .IN1(n6775), .IN2(n6100), .IN3(\FIFO[20][28] ), .IN4(n6104), 
        .Q(n3919) );
  AO22X1 U3848 ( .IN1(n6764), .IN2(n6101), .IN3(\FIFO[20][29] ), .IN4(n6104), 
        .Q(n3920) );
  AO22X1 U3849 ( .IN1(n6753), .IN2(n6100), .IN3(\FIFO[20][30] ), .IN4(n6104), 
        .Q(n3921) );
  AO22X1 U3850 ( .IN1(n6742), .IN2(n6099), .IN3(\FIFO[20][31] ), .IN4(n6104), 
        .Q(n3922) );
  AO21X1 U3851 ( .IN1(n357), .IN2(n261), .IN3(n7361), .Q(n368) );
  AO22X1 U3876 ( .IN1(n6819), .IN2(n369), .IN3(\FIFO[19][24] ), .IN4(n6098), 
        .Q(n3947) );
  AO22X1 U3877 ( .IN1(n6808), .IN2(n369), .IN3(\FIFO[19][25] ), .IN4(n6098), 
        .Q(n3948) );
  AO22X1 U3878 ( .IN1(n6797), .IN2(n369), .IN3(\FIFO[19][26] ), .IN4(n6098), 
        .Q(n3949) );
  AO22X1 U3879 ( .IN1(n6786), .IN2(n6095), .IN3(\FIFO[19][27] ), .IN4(n6098), 
        .Q(n3950) );
  AO22X1 U3880 ( .IN1(n6775), .IN2(n6094), .IN3(\FIFO[19][28] ), .IN4(n6098), 
        .Q(n3951) );
  AO22X1 U3881 ( .IN1(n6764), .IN2(n6095), .IN3(\FIFO[19][29] ), .IN4(n6098), 
        .Q(n3952) );
  AO22X1 U3882 ( .IN1(n6753), .IN2(n6094), .IN3(\FIFO[19][30] ), .IN4(n6098), 
        .Q(n3953) );
  AO22X1 U3883 ( .IN1(n6742), .IN2(n6093), .IN3(\FIFO[19][31] ), .IN4(n6098), 
        .Q(n3954) );
  AO21X1 U3884 ( .IN1(n357), .IN2(n263), .IN3(n7361), .Q(n369) );
  AO22X1 U3909 ( .IN1(n6819), .IN2(n370), .IN3(\FIFO[18][24] ), .IN4(n6092), 
        .Q(n3979) );
  AO22X1 U3910 ( .IN1(n6808), .IN2(n370), .IN3(\FIFO[18][25] ), .IN4(n6092), 
        .Q(n3980) );
  AO22X1 U3911 ( .IN1(n6797), .IN2(n370), .IN3(\FIFO[18][26] ), .IN4(n6092), 
        .Q(n3981) );
  AO22X1 U3912 ( .IN1(n6786), .IN2(n6089), .IN3(\FIFO[18][27] ), .IN4(n6092), 
        .Q(n3982) );
  AO22X1 U3913 ( .IN1(n6775), .IN2(n6089), .IN3(\FIFO[18][28] ), .IN4(n6092), 
        .Q(n3983) );
  AO22X1 U3914 ( .IN1(n6764), .IN2(n6088), .IN3(\FIFO[18][29] ), .IN4(n6092), 
        .Q(n3984) );
  AO22X1 U3915 ( .IN1(n6753), .IN2(n6087), .IN3(\FIFO[18][30] ), .IN4(n6092), 
        .Q(n3985) );
  AO22X1 U3916 ( .IN1(n6742), .IN2(n6088), .IN3(\FIFO[18][31] ), .IN4(n6092), 
        .Q(n3986) );
  AO21X1 U3917 ( .IN1(n357), .IN2(n265), .IN3(n7361), .Q(n370) );
  AO22X1 U3918 ( .IN1(n7089), .IN2(n6083), .IN3(\FIFO[17][0] ), .IN4(n6084), 
        .Q(n3987) );
  AO22X1 U3919 ( .IN1(n7072), .IN2(n6083), .IN3(\FIFO[17][1] ), .IN4(n6084), 
        .Q(n3988) );
  AO22X1 U3920 ( .IN1(n7061), .IN2(n6083), .IN3(\FIFO[17][2] ), .IN4(n6084), 
        .Q(n3989) );
  AO22X1 U3921 ( .IN1(n7050), .IN2(n6083), .IN3(\FIFO[17][3] ), .IN4(n6084), 
        .Q(n3990) );
  AO22X1 U3922 ( .IN1(n7039), .IN2(n6083), .IN3(\FIFO[17][4] ), .IN4(n6084), 
        .Q(n3991) );
  AO22X1 U3923 ( .IN1(n7028), .IN2(n6083), .IN3(\FIFO[17][5] ), .IN4(n6084), 
        .Q(n3992) );
  AO22X1 U3924 ( .IN1(n7017), .IN2(n6083), .IN3(\FIFO[17][6] ), .IN4(n6084), 
        .Q(n3993) );
  AO22X1 U3925 ( .IN1(n7006), .IN2(n6082), .IN3(\FIFO[17][7] ), .IN4(n6084), 
        .Q(n3994) );
  AO22X1 U3926 ( .IN1(n6995), .IN2(n6082), .IN3(\FIFO[17][8] ), .IN4(n6084), 
        .Q(n3995) );
  AO22X1 U3927 ( .IN1(n6984), .IN2(n6082), .IN3(\FIFO[17][9] ), .IN4(n6084), 
        .Q(n3996) );
  AO22X1 U3928 ( .IN1(n6973), .IN2(n6082), .IN3(\FIFO[17][10] ), .IN4(n6084), 
        .Q(n3997) );
  AO22X1 U3930 ( .IN1(n6951), .IN2(n6082), .IN3(\FIFO[17][12] ), .IN4(n6085), 
        .Q(n3999) );
  AO22X1 U3931 ( .IN1(n6940), .IN2(n6082), .IN3(\FIFO[17][13] ), .IN4(n6085), 
        .Q(n4000) );
  AO22X1 U3932 ( .IN1(n6929), .IN2(n6083), .IN3(\FIFO[17][14] ), .IN4(n6085), 
        .Q(n4001) );
  AO22X1 U3933 ( .IN1(n6918), .IN2(n6082), .IN3(\FIFO[17][15] ), .IN4(n6085), 
        .Q(n4002) );
  AO22X1 U3935 ( .IN1(n6896), .IN2(n6083), .IN3(\FIFO[17][17] ), .IN4(n6085), 
        .Q(n4004) );
  AO22X1 U3936 ( .IN1(n6885), .IN2(n6082), .IN3(\FIFO[17][18] ), .IN4(n6085), 
        .Q(n4005) );
  AO22X1 U3937 ( .IN1(n6874), .IN2(n6081), .IN3(\FIFO[17][19] ), .IN4(n6085), 
        .Q(n4006) );
  AO22X1 U3938 ( .IN1(n6863), .IN2(n6083), .IN3(\FIFO[17][20] ), .IN4(n6085), 
        .Q(n4007) );
  AO22X1 U3939 ( .IN1(n6852), .IN2(n6081), .IN3(\FIFO[17][21] ), .IN4(n6085), 
        .Q(n4008) );
  AO22X1 U3940 ( .IN1(n6841), .IN2(n6081), .IN3(\FIFO[17][22] ), .IN4(n6085), 
        .Q(n4009) );
  AO22X1 U3941 ( .IN1(n6830), .IN2(n6081), .IN3(\FIFO[17][23] ), .IN4(n6085), 
        .Q(n4010) );
  AO22X1 U3943 ( .IN1(n6808), .IN2(n6081), .IN3(\FIFO[17][25] ), .IN4(n6086), 
        .Q(n4012) );
  AO22X1 U3944 ( .IN1(n6797), .IN2(n6081), .IN3(\FIFO[17][26] ), .IN4(n6086), 
        .Q(n4013) );
  AO22X1 U3945 ( .IN1(n6786), .IN2(n6081), .IN3(\FIFO[17][27] ), .IN4(n6086), 
        .Q(n4014) );
  AO22X1 U3946 ( .IN1(n6775), .IN2(n6081), .IN3(\FIFO[17][28] ), .IN4(n6086), 
        .Q(n4015) );
  AO22X1 U3947 ( .IN1(n6764), .IN2(n6082), .IN3(\FIFO[17][29] ), .IN4(n6086), 
        .Q(n4016) );
  AO22X1 U3948 ( .IN1(n6753), .IN2(n6081), .IN3(\FIFO[17][30] ), .IN4(n6086), 
        .Q(n4017) );
  AO22X1 U3949 ( .IN1(n6742), .IN2(n6082), .IN3(\FIFO[17][31] ), .IN4(n6086), 
        .Q(n4018) );
  AO21X1 U3950 ( .IN1(n357), .IN2(n267), .IN3(n7361), .Q(n371) );
  AO22X1 U3951 ( .IN1(n7089), .IN2(n6077), .IN3(\FIFO[16][0] ), .IN4(n6078), 
        .Q(n4019) );
  AO22X1 U3952 ( .IN1(n7072), .IN2(n6076), .IN3(\FIFO[16][1] ), .IN4(n6078), 
        .Q(n4020) );
  AO22X1 U3953 ( .IN1(n7061), .IN2(n6075), .IN3(\FIFO[16][2] ), .IN4(n6078), 
        .Q(n4021) );
  AO22X1 U3954 ( .IN1(n7050), .IN2(n6077), .IN3(\FIFO[16][3] ), .IN4(n6078), 
        .Q(n4022) );
  AO22X1 U3955 ( .IN1(n7039), .IN2(n6076), .IN3(\FIFO[16][4] ), .IN4(n6078), 
        .Q(n4023) );
  AO22X1 U3957 ( .IN1(n7017), .IN2(n6077), .IN3(\FIFO[16][6] ), .IN4(n6078), 
        .Q(n4025) );
  AO22X1 U3958 ( .IN1(n7006), .IN2(n6077), .IN3(\FIFO[16][7] ), .IN4(n6078), 
        .Q(n4026) );
  AO22X1 U3959 ( .IN1(n6995), .IN2(n6077), .IN3(\FIFO[16][8] ), .IN4(n6078), 
        .Q(n4027) );
  AO22X1 U3960 ( .IN1(n6984), .IN2(n6077), .IN3(\FIFO[16][9] ), .IN4(n6078), 
        .Q(n4028) );
  AO22X1 U3961 ( .IN1(n6973), .IN2(n6077), .IN3(\FIFO[16][10] ), .IN4(n6078), 
        .Q(n4029) );
  AO22X1 U3962 ( .IN1(n6962), .IN2(n6077), .IN3(\FIFO[16][11] ), .IN4(n6078), 
        .Q(n4030) );
  AO22X1 U3963 ( .IN1(n6951), .IN2(n6077), .IN3(\FIFO[16][12] ), .IN4(n6079), 
        .Q(n4031) );
  AO22X1 U3964 ( .IN1(n6940), .IN2(n6077), .IN3(\FIFO[16][13] ), .IN4(n6079), 
        .Q(n4032) );
  AO22X1 U3965 ( .IN1(n6929), .IN2(n6076), .IN3(\FIFO[16][14] ), .IN4(n6079), 
        .Q(n4033) );
  AO22X1 U3966 ( .IN1(n6918), .IN2(n6076), .IN3(\FIFO[16][15] ), .IN4(n6079), 
        .Q(n4034) );
  AO22X1 U3967 ( .IN1(n6907), .IN2(n6076), .IN3(\FIFO[16][16] ), .IN4(n6079), 
        .Q(n4035) );
  AO22X1 U3969 ( .IN1(n6885), .IN2(n6076), .IN3(\FIFO[16][18] ), .IN4(n6079), 
        .Q(n4037) );
  AO22X1 U3970 ( .IN1(n6874), .IN2(n6076), .IN3(\FIFO[16][19] ), .IN4(n6079), 
        .Q(n4038) );
  AO22X1 U3971 ( .IN1(n6863), .IN2(n6076), .IN3(\FIFO[16][20] ), .IN4(n6079), 
        .Q(n4039) );
  AO22X1 U3972 ( .IN1(n6852), .IN2(n6075), .IN3(\FIFO[16][21] ), .IN4(n6079), 
        .Q(n4040) );
  AO22X1 U3973 ( .IN1(n6841), .IN2(n6075), .IN3(\FIFO[16][22] ), .IN4(n6079), 
        .Q(n4041) );
  AO22X1 U3974 ( .IN1(n6830), .IN2(n6075), .IN3(\FIFO[16][23] ), .IN4(n6079), 
        .Q(n4042) );
  AO22X1 U3975 ( .IN1(n6819), .IN2(n6075), .IN3(\FIFO[16][24] ), .IN4(n6080), 
        .Q(n4043) );
  AO22X1 U3977 ( .IN1(n6797), .IN2(n6075), .IN3(\FIFO[16][26] ), .IN4(n6080), 
        .Q(n4045) );
  AO22X1 U3978 ( .IN1(n6786), .IN2(n6075), .IN3(\FIFO[16][27] ), .IN4(n6080), 
        .Q(n4046) );
  AO22X1 U3979 ( .IN1(n6775), .IN2(n6075), .IN3(\FIFO[16][28] ), .IN4(n6080), 
        .Q(n4047) );
  AO22X1 U3980 ( .IN1(n6764), .IN2(n6076), .IN3(\FIFO[16][29] ), .IN4(n6080), 
        .Q(n4048) );
  AO22X1 U3981 ( .IN1(n6753), .IN2(n6075), .IN3(\FIFO[16][30] ), .IN4(n6080), 
        .Q(n4049) );
  AO22X1 U3982 ( .IN1(n6742), .IN2(n6076), .IN3(\FIFO[16][31] ), .IN4(n6080), 
        .Q(n4050) );
  AO21X1 U3983 ( .IN1(n357), .IN2(n269), .IN3(n7361), .Q(n372) );
  AO22X1 U4009 ( .IN1(n6819), .IN2(n373), .IN3(\FIFO[15][24] ), .IN4(n6074), 
        .Q(n4075) );
  AO22X1 U4010 ( .IN1(n6808), .IN2(n373), .IN3(\FIFO[15][25] ), .IN4(n6074), 
        .Q(n4076) );
  AO22X1 U4011 ( .IN1(n6797), .IN2(n373), .IN3(\FIFO[15][26] ), .IN4(n6074), 
        .Q(n4077) );
  AO22X1 U4012 ( .IN1(n6786), .IN2(n6071), .IN3(\FIFO[15][27] ), .IN4(n6074), 
        .Q(n4078) );
  AO22X1 U4013 ( .IN1(n6775), .IN2(n6070), .IN3(\FIFO[15][28] ), .IN4(n6074), 
        .Q(n4079) );
  AO22X1 U4014 ( .IN1(n6764), .IN2(n6071), .IN3(\FIFO[15][29] ), .IN4(n6074), 
        .Q(n4080) );
  AO22X1 U4015 ( .IN1(n6753), .IN2(n6070), .IN3(\FIFO[15][30] ), .IN4(n6074), 
        .Q(n4081) );
  AO22X1 U4016 ( .IN1(n6742), .IN2(n6069), .IN3(\FIFO[15][31] ), .IN4(n6074), 
        .Q(n4082) );
  AO22X1 U4043 ( .IN1(n6819), .IN2(n377), .IN3(\FIFO[14][24] ), .IN4(n6068), 
        .Q(n4107) );
  AO22X1 U4044 ( .IN1(n6808), .IN2(n377), .IN3(\FIFO[14][25] ), .IN4(n6068), 
        .Q(n4108) );
  AO22X1 U4045 ( .IN1(n6797), .IN2(n377), .IN3(\FIFO[14][26] ), .IN4(n6068), 
        .Q(n4109) );
  AO22X1 U4046 ( .IN1(n6786), .IN2(n6065), .IN3(\FIFO[14][27] ), .IN4(n6068), 
        .Q(n4110) );
  AO22X1 U4047 ( .IN1(n6775), .IN2(n6065), .IN3(\FIFO[14][28] ), .IN4(n6068), 
        .Q(n4111) );
  AO22X1 U4048 ( .IN1(n6764), .IN2(n6064), .IN3(\FIFO[14][29] ), .IN4(n6068), 
        .Q(n4112) );
  AO22X1 U4049 ( .IN1(n6753), .IN2(n6063), .IN3(\FIFO[14][30] ), .IN4(n6068), 
        .Q(n4113) );
  AO22X1 U4050 ( .IN1(n6742), .IN2(n6064), .IN3(\FIFO[14][31] ), .IN4(n6068), 
        .Q(n4114) );
  AO22X1 U4053 ( .IN1(n7089), .IN2(n6059), .IN3(\FIFO[13][0] ), .IN4(n6060), 
        .Q(n4115) );
  AO22X1 U4054 ( .IN1(n7072), .IN2(n6059), .IN3(\FIFO[13][1] ), .IN4(n6060), 
        .Q(n4116) );
  AO22X1 U4055 ( .IN1(n7061), .IN2(n6059), .IN3(\FIFO[13][2] ), .IN4(n6060), 
        .Q(n4117) );
  AO22X1 U4056 ( .IN1(n7050), .IN2(n6059), .IN3(\FIFO[13][3] ), .IN4(n6060), 
        .Q(n4118) );
  AO22X1 U4057 ( .IN1(n7039), .IN2(n6059), .IN3(\FIFO[13][4] ), .IN4(n6060), 
        .Q(n4119) );
  AO22X1 U4058 ( .IN1(n7028), .IN2(n6059), .IN3(\FIFO[13][5] ), .IN4(n6060), 
        .Q(n4120) );
  AO22X1 U4060 ( .IN1(n7006), .IN2(n6058), .IN3(\FIFO[13][7] ), .IN4(n6060), 
        .Q(n4122) );
  AO22X1 U4061 ( .IN1(n6995), .IN2(n6058), .IN3(\FIFO[13][8] ), .IN4(n6060), 
        .Q(n4123) );
  AO22X1 U4062 ( .IN1(n6984), .IN2(n6058), .IN3(\FIFO[13][9] ), .IN4(n6060), 
        .Q(n4124) );
  AO22X1 U4063 ( .IN1(n6973), .IN2(n6058), .IN3(\FIFO[13][10] ), .IN4(n6060), 
        .Q(n4125) );
  AO22X1 U4064 ( .IN1(n6962), .IN2(n6058), .IN3(\FIFO[13][11] ), .IN4(n6060), 
        .Q(n4126) );
  AO22X1 U4065 ( .IN1(n6951), .IN2(n6058), .IN3(\FIFO[13][12] ), .IN4(n6061), 
        .Q(n4127) );
  AO22X1 U4066 ( .IN1(n6940), .IN2(n6058), .IN3(\FIFO[13][13] ), .IN4(n6061), 
        .Q(n4128) );
  AO22X1 U4067 ( .IN1(n6929), .IN2(n6059), .IN3(\FIFO[13][14] ), .IN4(n6061), 
        .Q(n4129) );
  AO22X1 U4068 ( .IN1(n6918), .IN2(n6058), .IN3(\FIFO[13][15] ), .IN4(n6061), 
        .Q(n4130) );
  AO22X1 U4069 ( .IN1(n6907), .IN2(n6057), .IN3(\FIFO[13][16] ), .IN4(n6061), 
        .Q(n4131) );
  AO22X1 U4070 ( .IN1(n6896), .IN2(n6059), .IN3(\FIFO[13][17] ), .IN4(n6061), 
        .Q(n4132) );
  AO22X1 U4072 ( .IN1(n6874), .IN2(n6057), .IN3(\FIFO[13][19] ), .IN4(n6061), 
        .Q(n4134) );
  AO22X1 U4073 ( .IN1(n6863), .IN2(n6059), .IN3(\FIFO[13][20] ), .IN4(n6061), 
        .Q(n4135) );
  AO22X1 U4074 ( .IN1(n6852), .IN2(n6057), .IN3(\FIFO[13][21] ), .IN4(n6061), 
        .Q(n4136) );
  AO22X1 U4075 ( .IN1(n6841), .IN2(n6057), .IN3(\FIFO[13][22] ), .IN4(n6061), 
        .Q(n4137) );
  AO22X1 U4076 ( .IN1(n6830), .IN2(n6057), .IN3(\FIFO[13][23] ), .IN4(n6061), 
        .Q(n4138) );
  AO22X1 U4077 ( .IN1(n6819), .IN2(n6057), .IN3(\FIFO[13][24] ), .IN4(n6062), 
        .Q(n4139) );
  AO22X1 U4078 ( .IN1(n6808), .IN2(n6057), .IN3(\FIFO[13][25] ), .IN4(n6062), 
        .Q(n4140) );
  AO22X1 U4080 ( .IN1(n6786), .IN2(n6057), .IN3(\FIFO[13][27] ), .IN4(n6062), 
        .Q(n4142) );
  AO22X1 U4081 ( .IN1(n6775), .IN2(n6057), .IN3(\FIFO[13][28] ), .IN4(n6062), 
        .Q(n4143) );
  AO22X1 U4082 ( .IN1(n6764), .IN2(n6058), .IN3(\FIFO[13][29] ), .IN4(n6062), 
        .Q(n4144) );
  AO22X1 U4083 ( .IN1(n6753), .IN2(n6057), .IN3(\FIFO[13][30] ), .IN4(n6062), 
        .Q(n4145) );
  AO22X1 U4084 ( .IN1(n6742), .IN2(n6058), .IN3(\FIFO[13][31] ), .IN4(n6062), 
        .Q(n4146) );
  AO21X1 U4085 ( .IN1(n374), .IN2(n243), .IN3(n7361), .Q(n379) );
  AND2X1 U4086 ( .IN1(n380), .IN2(n375), .Q(n243) );
  AO22X1 U4087 ( .IN1(n7089), .IN2(n6053), .IN3(\FIFO[12][0] ), .IN4(n6054), 
        .Q(n4147) );
  AO22X1 U4088 ( .IN1(n7072), .IN2(n6052), .IN3(\FIFO[12][1] ), .IN4(n6054), 
        .Q(n4148) );
  AO22X1 U4089 ( .IN1(n7061), .IN2(n6051), .IN3(\FIFO[12][2] ), .IN4(n6054), 
        .Q(n4149) );
  AO22X1 U4090 ( .IN1(n7050), .IN2(n6053), .IN3(\FIFO[12][3] ), .IN4(n6054), 
        .Q(n4150) );
  AO22X1 U4091 ( .IN1(n7039), .IN2(n6052), .IN3(\FIFO[12][4] ), .IN4(n6054), 
        .Q(n4151) );
  AO22X1 U4092 ( .IN1(n7028), .IN2(n6051), .IN3(\FIFO[12][5] ), .IN4(n6054), 
        .Q(n4152) );
  AO22X1 U4093 ( .IN1(n7017), .IN2(n6053), .IN3(\FIFO[12][6] ), .IN4(n6054), 
        .Q(n4153) );
  AO22X1 U4095 ( .IN1(n6995), .IN2(n6053), .IN3(\FIFO[12][8] ), .IN4(n6054), 
        .Q(n4155) );
  AO22X1 U4096 ( .IN1(n6984), .IN2(n6053), .IN3(\FIFO[12][9] ), .IN4(n6054), 
        .Q(n4156) );
  AO22X1 U4097 ( .IN1(n6973), .IN2(n6053), .IN3(\FIFO[12][10] ), .IN4(n6054), 
        .Q(n4157) );
  AO22X1 U4098 ( .IN1(n6962), .IN2(n6053), .IN3(\FIFO[12][11] ), .IN4(n6054), 
        .Q(n4158) );
  AO22X1 U4099 ( .IN1(n6951), .IN2(n6053), .IN3(\FIFO[12][12] ), .IN4(n6055), 
        .Q(n4159) );
  AO22X1 U4100 ( .IN1(n6940), .IN2(n6053), .IN3(\FIFO[12][13] ), .IN4(n6055), 
        .Q(n4160) );
  AO22X1 U4101 ( .IN1(n6929), .IN2(n6052), .IN3(\FIFO[12][14] ), .IN4(n6055), 
        .Q(n4161) );
  AO22X1 U4102 ( .IN1(n6918), .IN2(n6052), .IN3(\FIFO[12][15] ), .IN4(n6055), 
        .Q(n4162) );
  AO22X1 U4103 ( .IN1(n6907), .IN2(n6052), .IN3(\FIFO[12][16] ), .IN4(n6055), 
        .Q(n4163) );
  AO22X1 U4104 ( .IN1(n6896), .IN2(n6052), .IN3(\FIFO[12][17] ), .IN4(n6055), 
        .Q(n4164) );
  AO22X1 U4105 ( .IN1(n6885), .IN2(n6052), .IN3(\FIFO[12][18] ), .IN4(n6055), 
        .Q(n4165) );
  AO22X1 U4107 ( .IN1(n6863), .IN2(n6052), .IN3(\FIFO[12][20] ), .IN4(n6055), 
        .Q(n4167) );
  AO22X1 U4108 ( .IN1(n6852), .IN2(n6051), .IN3(\FIFO[12][21] ), .IN4(n6055), 
        .Q(n4168) );
  AO22X1 U4109 ( .IN1(n6841), .IN2(n6051), .IN3(\FIFO[12][22] ), .IN4(n6055), 
        .Q(n4169) );
  AO22X1 U4110 ( .IN1(n6830), .IN2(n6051), .IN3(\FIFO[12][23] ), .IN4(n6055), 
        .Q(n4170) );
  AO22X1 U4111 ( .IN1(n6819), .IN2(n6051), .IN3(\FIFO[12][24] ), .IN4(n6056), 
        .Q(n4171) );
  AO22X1 U4112 ( .IN1(n6808), .IN2(n6051), .IN3(\FIFO[12][25] ), .IN4(n6056), 
        .Q(n4172) );
  AO22X1 U4113 ( .IN1(n6797), .IN2(n6051), .IN3(\FIFO[12][26] ), .IN4(n6056), 
        .Q(n4173) );
  AO22X1 U4115 ( .IN1(n6775), .IN2(n6051), .IN3(\FIFO[12][28] ), .IN4(n6056), 
        .Q(n4175) );
  AO22X1 U4116 ( .IN1(n6764), .IN2(n6052), .IN3(\FIFO[12][29] ), .IN4(n6056), 
        .Q(n4176) );
  AO22X1 U4117 ( .IN1(n6753), .IN2(n6051), .IN3(\FIFO[12][30] ), .IN4(n6056), 
        .Q(n4177) );
  AO22X1 U4118 ( .IN1(n6742), .IN2(n6052), .IN3(\FIFO[12][31] ), .IN4(n6056), 
        .Q(n4178) );
  AO21X1 U4119 ( .IN1(n374), .IN2(n245), .IN3(n7361), .Q(n381) );
  AND2X1 U4120 ( .IN1(n382), .IN2(n375), .Q(n245) );
  AO22X1 U4145 ( .IN1(n6818), .IN2(n383), .IN3(\FIFO[11][24] ), .IN4(n6050), 
        .Q(n4203) );
  AO22X1 U4146 ( .IN1(n6807), .IN2(n383), .IN3(\FIFO[11][25] ), .IN4(n6050), 
        .Q(n4204) );
  AO22X1 U4147 ( .IN1(n6796), .IN2(n383), .IN3(\FIFO[11][26] ), .IN4(n6050), 
        .Q(n4205) );
  AO22X1 U4148 ( .IN1(n6785), .IN2(n6047), .IN3(\FIFO[11][27] ), .IN4(n6050), 
        .Q(n4206) );
  AO22X1 U4149 ( .IN1(n6774), .IN2(n6046), .IN3(\FIFO[11][28] ), .IN4(n6050), 
        .Q(n4207) );
  AO22X1 U4150 ( .IN1(n6763), .IN2(n6047), .IN3(\FIFO[11][29] ), .IN4(n6050), 
        .Q(n4208) );
  AO22X1 U4151 ( .IN1(n6752), .IN2(n6046), .IN3(\FIFO[11][30] ), .IN4(n6050), 
        .Q(n4209) );
  AO22X1 U4152 ( .IN1(n6741), .IN2(n6045), .IN3(\FIFO[11][31] ), .IN4(n6050), 
        .Q(n4210) );
  AO22X1 U4179 ( .IN1(n6818), .IN2(n385), .IN3(\FIFO[10][24] ), .IN4(n6044), 
        .Q(n4235) );
  AO22X1 U4180 ( .IN1(n6807), .IN2(n385), .IN3(\FIFO[10][25] ), .IN4(n6044), 
        .Q(n4236) );
  AO22X1 U4181 ( .IN1(n6796), .IN2(n385), .IN3(\FIFO[10][26] ), .IN4(n6044), 
        .Q(n4237) );
  AO22X1 U4182 ( .IN1(n6785), .IN2(n6041), .IN3(\FIFO[10][27] ), .IN4(n6044), 
        .Q(n4238) );
  AO22X1 U4183 ( .IN1(n6774), .IN2(n6040), .IN3(\FIFO[10][28] ), .IN4(n6044), 
        .Q(n4239) );
  AO22X1 U4184 ( .IN1(n6763), .IN2(n6041), .IN3(\FIFO[10][29] ), .IN4(n6044), 
        .Q(n4240) );
  AO22X1 U4185 ( .IN1(n6752), .IN2(n6040), .IN3(\FIFO[10][30] ), .IN4(n6044), 
        .Q(n4241) );
  AO22X1 U4186 ( .IN1(n6741), .IN2(n6039), .IN3(\FIFO[10][31] ), .IN4(n6044), 
        .Q(n4242) );
  AO22X1 U4189 ( .IN1(n7088), .IN2(n6035), .IN3(\FIFO[9][0] ), .IN4(n6036), 
        .Q(n4243) );
  AO22X1 U4190 ( .IN1(n7071), .IN2(n6035), .IN3(\FIFO[9][1] ), .IN4(n6036), 
        .Q(n4244) );
  AO22X1 U4191 ( .IN1(n7060), .IN2(n6035), .IN3(\FIFO[9][2] ), .IN4(n6036), 
        .Q(n4245) );
  AO22X1 U4192 ( .IN1(n7049), .IN2(n6035), .IN3(\FIFO[9][3] ), .IN4(n6036), 
        .Q(n4246) );
  AO22X1 U4193 ( .IN1(n7038), .IN2(n6035), .IN3(\FIFO[9][4] ), .IN4(n6036), 
        .Q(n4247) );
  AO22X1 U4194 ( .IN1(n7027), .IN2(n6035), .IN3(\FIFO[9][5] ), .IN4(n6036), 
        .Q(n4248) );
  AO22X1 U4195 ( .IN1(n7016), .IN2(n6035), .IN3(\FIFO[9][6] ), .IN4(n6036), 
        .Q(n4249) );
  AO22X1 U4197 ( .IN1(n6994), .IN2(n6034), .IN3(\FIFO[9][8] ), .IN4(n6036), 
        .Q(n4251) );
  AO22X1 U4198 ( .IN1(n6983), .IN2(n6034), .IN3(\FIFO[9][9] ), .IN4(n6036), 
        .Q(n4252) );
  AO22X1 U4199 ( .IN1(n6972), .IN2(n6034), .IN3(\FIFO[9][10] ), .IN4(n6036), 
        .Q(n4253) );
  AO22X1 U4200 ( .IN1(n6961), .IN2(n6034), .IN3(\FIFO[9][11] ), .IN4(n6036), 
        .Q(n4254) );
  AO22X1 U4201 ( .IN1(n6950), .IN2(n6034), .IN3(\FIFO[9][12] ), .IN4(n6037), 
        .Q(n4255) );
  AO22X1 U4202 ( .IN1(n6939), .IN2(n6034), .IN3(\FIFO[9][13] ), .IN4(n6037), 
        .Q(n4256) );
  AO22X1 U4203 ( .IN1(n6928), .IN2(n6033), .IN3(\FIFO[9][14] ), .IN4(n6037), 
        .Q(n4257) );
  AO22X1 U4204 ( .IN1(n6917), .IN2(n6033), .IN3(\FIFO[9][15] ), .IN4(n6037), 
        .Q(n4258) );
  AO22X1 U4205 ( .IN1(n6906), .IN2(n6033), .IN3(\FIFO[9][16] ), .IN4(n6037), 
        .Q(n4259) );
  AO22X1 U4206 ( .IN1(n6895), .IN2(n6033), .IN3(\FIFO[9][17] ), .IN4(n6037), 
        .Q(n4260) );
  AO22X1 U4208 ( .IN1(n6873), .IN2(n6033), .IN3(\FIFO[9][19] ), .IN4(n6037), 
        .Q(n4262) );
  AO22X1 U4209 ( .IN1(n6862), .IN2(n6033), .IN3(\FIFO[9][20] ), .IN4(n6037), 
        .Q(n4263) );
  AO22X1 U4210 ( .IN1(n6851), .IN2(n6035), .IN3(\FIFO[9][21] ), .IN4(n6037), 
        .Q(n4264) );
  AO22X1 U4211 ( .IN1(n6840), .IN2(n6034), .IN3(\FIFO[9][22] ), .IN4(n6037), 
        .Q(n4265) );
  AO22X1 U4212 ( .IN1(n6829), .IN2(n6033), .IN3(\FIFO[9][23] ), .IN4(n6037), 
        .Q(n4266) );
  AO22X1 U4213 ( .IN1(n6818), .IN2(n386), .IN3(\FIFO[9][24] ), .IN4(n6038), 
        .Q(n4267) );
  AO22X1 U4214 ( .IN1(n6807), .IN2(n386), .IN3(\FIFO[9][25] ), .IN4(n6038), 
        .Q(n4268) );
  AO22X1 U4215 ( .IN1(n6796), .IN2(n386), .IN3(\FIFO[9][26] ), .IN4(n6038), 
        .Q(n4269) );
  AO22X1 U4216 ( .IN1(n6785), .IN2(n6035), .IN3(\FIFO[9][27] ), .IN4(n6038), 
        .Q(n4270) );
  AO22X1 U4217 ( .IN1(n6774), .IN2(n6035), .IN3(\FIFO[9][28] ), .IN4(n6038), 
        .Q(n4271) );
  AO22X1 U4218 ( .IN1(n6763), .IN2(n6034), .IN3(\FIFO[9][29] ), .IN4(n6038), 
        .Q(n4272) );
  AO22X1 U4219 ( .IN1(n6752), .IN2(n6033), .IN3(\FIFO[9][30] ), .IN4(n6038), 
        .Q(n4273) );
  AO22X1 U4220 ( .IN1(n6741), .IN2(n6034), .IN3(\FIFO[9][31] ), .IN4(n6038), 
        .Q(n4274) );
  AO22X1 U4223 ( .IN1(n7088), .IN2(n6029), .IN3(\FIFO[8][0] ), .IN4(n6030), 
        .Q(n4275) );
  AO22X1 U4224 ( .IN1(n7071), .IN2(n6029), .IN3(\FIFO[8][1] ), .IN4(n6030), 
        .Q(n4276) );
  AO22X1 U4225 ( .IN1(n7060), .IN2(n6029), .IN3(\FIFO[8][2] ), .IN4(n6030), 
        .Q(n4277) );
  AO22X1 U4226 ( .IN1(n7049), .IN2(n6029), .IN3(\FIFO[8][3] ), .IN4(n6030), 
        .Q(n4278) );
  AO22X1 U4227 ( .IN1(n7038), .IN2(n6029), .IN3(\FIFO[8][4] ), .IN4(n6030), 
        .Q(n4279) );
  AO22X1 U4228 ( .IN1(n7027), .IN2(n6029), .IN3(\FIFO[8][5] ), .IN4(n6030), 
        .Q(n4280) );
  AO22X1 U4229 ( .IN1(n7016), .IN2(n6029), .IN3(\FIFO[8][6] ), .IN4(n6030), 
        .Q(n4281) );
  AO22X1 U4230 ( .IN1(n7005), .IN2(n6028), .IN3(\FIFO[8][7] ), .IN4(n6030), 
        .Q(n4282) );
  AO22X1 U4231 ( .IN1(n6994), .IN2(n6028), .IN3(\FIFO[8][8] ), .IN4(n6030), 
        .Q(n4283) );
  AO22X1 U4232 ( .IN1(n6983), .IN2(n6028), .IN3(\FIFO[8][9] ), .IN4(n6030), 
        .Q(n4284) );
  AO22X1 U4233 ( .IN1(n6972), .IN2(n6028), .IN3(\FIFO[8][10] ), .IN4(n6030), 
        .Q(n4285) );
  AO22X1 U4234 ( .IN1(n6961), .IN2(n6028), .IN3(\FIFO[8][11] ), .IN4(n6030), 
        .Q(n4286) );
  AO22X1 U4235 ( .IN1(n6950), .IN2(n6028), .IN3(\FIFO[8][12] ), .IN4(n6031), 
        .Q(n4287) );
  AO22X1 U4237 ( .IN1(n6928), .IN2(n6029), .IN3(\FIFO[8][14] ), .IN4(n6031), 
        .Q(n4289) );
  AO22X1 U4238 ( .IN1(n6917), .IN2(n6028), .IN3(\FIFO[8][15] ), .IN4(n6031), 
        .Q(n4290) );
  AO22X1 U4239 ( .IN1(n6906), .IN2(n6027), .IN3(\FIFO[8][16] ), .IN4(n6031), 
        .Q(n4291) );
  AO22X1 U4240 ( .IN1(n6895), .IN2(n6029), .IN3(\FIFO[8][17] ), .IN4(n6031), 
        .Q(n4292) );
  AO22X1 U4241 ( .IN1(n6884), .IN2(n6028), .IN3(\FIFO[8][18] ), .IN4(n6031), 
        .Q(n4293) );
  AO22X1 U4242 ( .IN1(n6873), .IN2(n6027), .IN3(\FIFO[8][19] ), .IN4(n6031), 
        .Q(n4294) );
  AO22X1 U4244 ( .IN1(n6851), .IN2(n6027), .IN3(\FIFO[8][21] ), .IN4(n6031), 
        .Q(n4296) );
  AO22X1 U4245 ( .IN1(n6840), .IN2(n6027), .IN3(\FIFO[8][22] ), .IN4(n6031), 
        .Q(n4297) );
  AO22X1 U4246 ( .IN1(n6829), .IN2(n6027), .IN3(\FIFO[8][23] ), .IN4(n6031), 
        .Q(n4298) );
  AO22X1 U4247 ( .IN1(n6818), .IN2(n6027), .IN3(\FIFO[8][24] ), .IN4(n6032), 
        .Q(n4299) );
  AO22X1 U4248 ( .IN1(n6807), .IN2(n6027), .IN3(\FIFO[8][25] ), .IN4(n6032), 
        .Q(n4300) );
  AO22X1 U4249 ( .IN1(n6796), .IN2(n6027), .IN3(\FIFO[8][26] ), .IN4(n6032), 
        .Q(n4301) );
  AO22X1 U4250 ( .IN1(n6785), .IN2(n6027), .IN3(\FIFO[8][27] ), .IN4(n6032), 
        .Q(n4302) );
  AO22X1 U4252 ( .IN1(n6763), .IN2(n6028), .IN3(\FIFO[8][29] ), .IN4(n6032), 
        .Q(n4304) );
  AO22X1 U4253 ( .IN1(n6752), .IN2(n6027), .IN3(\FIFO[8][30] ), .IN4(n6032), 
        .Q(n4305) );
  AO22X1 U4254 ( .IN1(n6741), .IN2(n6028), .IN3(\FIFO[8][31] ), .IN4(n6032), 
        .Q(n4306) );
  AO21X1 U4255 ( .IN1(n374), .IN2(n253), .IN3(n7361), .Q(n387) );
  AND2X1 U4256 ( .IN1(n384), .IN2(n382), .Q(n253) );
  AO22X1 U4281 ( .IN1(n6818), .IN2(n6021), .IN3(\FIFO[7][24] ), .IN4(n6026), 
        .Q(n4331) );
  AO22X1 U4282 ( .IN1(n6807), .IN2(n6021), .IN3(\FIFO[7][25] ), .IN4(n6026), 
        .Q(n4332) );
  AO22X1 U4283 ( .IN1(n6796), .IN2(n6021), .IN3(\FIFO[7][26] ), .IN4(n6026), 
        .Q(n4333) );
  AO22X1 U4284 ( .IN1(n6785), .IN2(n6021), .IN3(\FIFO[7][27] ), .IN4(n6026), 
        .Q(n4334) );
  AO22X1 U4285 ( .IN1(n6774), .IN2(n6021), .IN3(\FIFO[7][28] ), .IN4(n6026), 
        .Q(n4335) );
  AO22X1 U4287 ( .IN1(n6752), .IN2(n6021), .IN3(\FIFO[7][30] ), .IN4(n6026), 
        .Q(n4337) );
  AO22X1 U4288 ( .IN1(n6741), .IN2(n6022), .IN3(\FIFO[7][31] ), .IN4(n6026), 
        .Q(n4338) );
  AO21X1 U4289 ( .IN1(n374), .IN2(n255), .IN3(n7361), .Q(n388) );
  AND2X1 U4290 ( .IN1(n389), .IN2(n376), .Q(n255) );
  AO22X1 U4315 ( .IN1(n6818), .IN2(n390), .IN3(\FIFO[6][24] ), .IN4(n6020), 
        .Q(n4363) );
  AO22X1 U4316 ( .IN1(n6807), .IN2(n390), .IN3(\FIFO[6][25] ), .IN4(n6020), 
        .Q(n4364) );
  AO22X1 U4317 ( .IN1(n6796), .IN2(n390), .IN3(\FIFO[6][26] ), .IN4(n6020), 
        .Q(n4365) );
  AO22X1 U4318 ( .IN1(n6785), .IN2(n6017), .IN3(\FIFO[6][27] ), .IN4(n6020), 
        .Q(n4366) );
  AO22X1 U4319 ( .IN1(n6774), .IN2(n6016), .IN3(\FIFO[6][28] ), .IN4(n6020), 
        .Q(n4367) );
  AO22X1 U4320 ( .IN1(n6763), .IN2(n6017), .IN3(\FIFO[6][29] ), .IN4(n6020), 
        .Q(n4368) );
  AO22X1 U4321 ( .IN1(n6752), .IN2(n6016), .IN3(\FIFO[6][30] ), .IN4(n6020), 
        .Q(n4369) );
  AO22X1 U4322 ( .IN1(n6741), .IN2(n6015), .IN3(\FIFO[6][31] ), .IN4(n6020), 
        .Q(n4370) );
  AO22X1 U4325 ( .IN1(n7088), .IN2(n6011), .IN3(\FIFO[5][0] ), .IN4(n6012), 
        .Q(n4371) );
  AO22X1 U4326 ( .IN1(n7071), .IN2(n6011), .IN3(\FIFO[5][1] ), .IN4(n6012), 
        .Q(n4372) );
  AO22X1 U4327 ( .IN1(n7060), .IN2(n6011), .IN3(\FIFO[5][2] ), .IN4(n6012), 
        .Q(n4373) );
  AO22X1 U4328 ( .IN1(n7049), .IN2(n6011), .IN3(\FIFO[5][3] ), .IN4(n6012), 
        .Q(n4374) );
  AO22X1 U4329 ( .IN1(n7038), .IN2(n6011), .IN3(\FIFO[5][4] ), .IN4(n6012), 
        .Q(n4375) );
  AO22X1 U4330 ( .IN1(n7027), .IN2(n6011), .IN3(\FIFO[5][5] ), .IN4(n6012), 
        .Q(n4376) );
  AO22X1 U4331 ( .IN1(n7016), .IN2(n6011), .IN3(\FIFO[5][6] ), .IN4(n6012), 
        .Q(n4377) );
  AO22X1 U4332 ( .IN1(n7005), .IN2(n6010), .IN3(\FIFO[5][7] ), .IN4(n6012), 
        .Q(n4378) );
  AO22X1 U4333 ( .IN1(n6994), .IN2(n6010), .IN3(\FIFO[5][8] ), .IN4(n6012), 
        .Q(n4379) );
  AO22X1 U4335 ( .IN1(n6972), .IN2(n6010), .IN3(\FIFO[5][10] ), .IN4(n6012), 
        .Q(n4381) );
  AO22X1 U4336 ( .IN1(n6961), .IN2(n6010), .IN3(\FIFO[5][11] ), .IN4(n6012), 
        .Q(n4382) );
  AO22X1 U4337 ( .IN1(n6950), .IN2(n6010), .IN3(\FIFO[5][12] ), .IN4(n6013), 
        .Q(n4383) );
  AO22X1 U4338 ( .IN1(n6939), .IN2(n6010), .IN3(\FIFO[5][13] ), .IN4(n6013), 
        .Q(n4384) );
  AO22X1 U4339 ( .IN1(n6928), .IN2(n6009), .IN3(\FIFO[5][14] ), .IN4(n6013), 
        .Q(n4385) );
  AO22X1 U4340 ( .IN1(n6917), .IN2(n6009), .IN3(\FIFO[5][15] ), .IN4(n6013), 
        .Q(n4386) );
  AO22X1 U4341 ( .IN1(n6906), .IN2(n6009), .IN3(\FIFO[5][16] ), .IN4(n6013), 
        .Q(n4387) );
  AO22X1 U4342 ( .IN1(n6895), .IN2(n6009), .IN3(\FIFO[5][17] ), .IN4(n6013), 
        .Q(n4388) );
  AO22X1 U4343 ( .IN1(n6884), .IN2(n6009), .IN3(\FIFO[5][18] ), .IN4(n6013), 
        .Q(n4389) );
  AO22X1 U4344 ( .IN1(n6873), .IN2(n6009), .IN3(\FIFO[5][19] ), .IN4(n6013), 
        .Q(n4390) );
  AO22X1 U4346 ( .IN1(n6851), .IN2(n6011), .IN3(\FIFO[5][21] ), .IN4(n6013), 
        .Q(n4392) );
  AO22X1 U4347 ( .IN1(n6840), .IN2(n6010), .IN3(\FIFO[5][22] ), .IN4(n6013), 
        .Q(n4393) );
  AO22X1 U4348 ( .IN1(n6829), .IN2(n6009), .IN3(\FIFO[5][23] ), .IN4(n6013), 
        .Q(n4394) );
  AO22X1 U4349 ( .IN1(n6818), .IN2(n391), .IN3(\FIFO[5][24] ), .IN4(n6014), 
        .Q(n4395) );
  AO22X1 U4350 ( .IN1(n6807), .IN2(n391), .IN3(\FIFO[5][25] ), .IN4(n6014), 
        .Q(n4396) );
  AO22X1 U4351 ( .IN1(n6796), .IN2(n391), .IN3(\FIFO[5][26] ), .IN4(n6014), 
        .Q(n4397) );
  AO22X1 U4352 ( .IN1(n6785), .IN2(n6011), .IN3(\FIFO[5][27] ), .IN4(n6014), 
        .Q(n4398) );
  AO22X1 U4353 ( .IN1(n6774), .IN2(n6010), .IN3(\FIFO[5][28] ), .IN4(n6014), 
        .Q(n4399) );
  AO22X1 U4354 ( .IN1(n6763), .IN2(n6011), .IN3(\FIFO[5][29] ), .IN4(n6014), 
        .Q(n4400) );
  AO22X1 U4355 ( .IN1(n6752), .IN2(n6010), .IN3(\FIFO[5][30] ), .IN4(n6014), 
        .Q(n4401) );
  AO22X1 U4356 ( .IN1(n6741), .IN2(n6009), .IN3(\FIFO[5][31] ), .IN4(n6014), 
        .Q(n4402) );
  AO22X1 U4359 ( .IN1(n7088), .IN2(n6005), .IN3(\FIFO[4][0] ), .IN4(n6006), 
        .Q(n4403) );
  AO22X1 U4360 ( .IN1(n7071), .IN2(n6005), .IN3(\FIFO[4][1] ), .IN4(n6006), 
        .Q(n4404) );
  AO22X1 U4361 ( .IN1(n7060), .IN2(n6005), .IN3(\FIFO[4][2] ), .IN4(n6006), 
        .Q(n4405) );
  AO22X1 U4362 ( .IN1(n7049), .IN2(n6005), .IN3(\FIFO[4][3] ), .IN4(n6006), 
        .Q(n4406) );
  AO22X1 U4363 ( .IN1(n7038), .IN2(n6005), .IN3(\FIFO[4][4] ), .IN4(n6006), 
        .Q(n4407) );
  AO22X1 U4364 ( .IN1(n7027), .IN2(n6005), .IN3(\FIFO[4][5] ), .IN4(n6006), 
        .Q(n4408) );
  AO22X1 U4365 ( .IN1(n7016), .IN2(n6005), .IN3(\FIFO[4][6] ), .IN4(n6006), 
        .Q(n4409) );
  AO22X1 U4366 ( .IN1(n7005), .IN2(n6004), .IN3(\FIFO[4][7] ), .IN4(n6006), 
        .Q(n4410) );
  AO22X1 U4367 ( .IN1(n6994), .IN2(n6004), .IN3(\FIFO[4][8] ), .IN4(n6006), 
        .Q(n4411) );
  AO22X1 U4368 ( .IN1(n6983), .IN2(n6004), .IN3(\FIFO[4][9] ), .IN4(n6006), 
        .Q(n4412) );
  AO22X1 U4370 ( .IN1(n6961), .IN2(n6004), .IN3(\FIFO[4][11] ), .IN4(n6006), 
        .Q(n4414) );
  AO22X1 U4371 ( .IN1(n6950), .IN2(n6004), .IN3(\FIFO[4][12] ), .IN4(n6007), 
        .Q(n4415) );
  AO22X1 U4372 ( .IN1(n6939), .IN2(n6004), .IN3(\FIFO[4][13] ), .IN4(n6007), 
        .Q(n4416) );
  AO22X1 U4373 ( .IN1(n6928), .IN2(n6003), .IN3(\FIFO[4][14] ), .IN4(n6007), 
        .Q(n4417) );
  AO22X1 U4374 ( .IN1(n6917), .IN2(n6003), .IN3(\FIFO[4][15] ), .IN4(n6007), 
        .Q(n4418) );
  AO22X1 U4375 ( .IN1(n6906), .IN2(n6003), .IN3(\FIFO[4][16] ), .IN4(n6007), 
        .Q(n4419) );
  AO22X1 U4376 ( .IN1(n6895), .IN2(n6003), .IN3(\FIFO[4][17] ), .IN4(n6007), 
        .Q(n4420) );
  AO22X1 U4377 ( .IN1(n6884), .IN2(n6003), .IN3(\FIFO[4][18] ), .IN4(n6007), 
        .Q(n4421) );
  AO22X1 U4378 ( .IN1(n6873), .IN2(n6003), .IN3(\FIFO[4][19] ), .IN4(n6007), 
        .Q(n4422) );
  AO22X1 U4379 ( .IN1(n6862), .IN2(n6003), .IN3(\FIFO[4][20] ), .IN4(n6007), 
        .Q(n4423) );
  AO22X1 U4381 ( .IN1(n6840), .IN2(n6004), .IN3(\FIFO[4][22] ), .IN4(n6007), 
        .Q(n4425) );
  AO22X1 U4382 ( .IN1(n6829), .IN2(n6003), .IN3(\FIFO[4][23] ), .IN4(n6007), 
        .Q(n4426) );
  AO22X1 U4383 ( .IN1(n6818), .IN2(n392), .IN3(\FIFO[4][24] ), .IN4(n6008), 
        .Q(n4427) );
  AO22X1 U4384 ( .IN1(n6807), .IN2(n392), .IN3(\FIFO[4][25] ), .IN4(n6008), 
        .Q(n4428) );
  AO22X1 U4385 ( .IN1(n6796), .IN2(n392), .IN3(\FIFO[4][26] ), .IN4(n6008), 
        .Q(n4429) );
  AO22X1 U4386 ( .IN1(n6785), .IN2(n6005), .IN3(\FIFO[4][27] ), .IN4(n6008), 
        .Q(n4430) );
  AO22X1 U4387 ( .IN1(n6774), .IN2(n6005), .IN3(\FIFO[4][28] ), .IN4(n6008), 
        .Q(n4431) );
  AO22X1 U4388 ( .IN1(n6763), .IN2(n6004), .IN3(\FIFO[4][29] ), .IN4(n6008), 
        .Q(n4432) );
  AO22X1 U4389 ( .IN1(n6752), .IN2(n6003), .IN3(\FIFO[4][30] ), .IN4(n6008), 
        .Q(n4433) );
  AO22X1 U4390 ( .IN1(n6741), .IN2(n6004), .IN3(\FIFO[4][31] ), .IN4(n6008), 
        .Q(n4434) );
  AO21X1 U4391 ( .IN1(n374), .IN2(n261), .IN3(n7361), .Q(n392) );
  AND2X1 U4392 ( .IN1(n389), .IN2(n382), .Q(n261) );
  AO22X1 U4417 ( .IN1(n6818), .IN2(n5997), .IN3(\FIFO[3][24] ), .IN4(n6002), 
        .Q(n4459) );
  AO22X1 U4418 ( .IN1(n6807), .IN2(n5997), .IN3(\FIFO[3][25] ), .IN4(n6002), 
        .Q(n4460) );
  AO22X1 U4419 ( .IN1(n6796), .IN2(n5997), .IN3(\FIFO[3][26] ), .IN4(n6002), 
        .Q(n4461) );
  AO22X1 U4420 ( .IN1(n6785), .IN2(n5997), .IN3(\FIFO[3][27] ), .IN4(n6002), 
        .Q(n4462) );
  AO22X1 U4421 ( .IN1(n6774), .IN2(n5997), .IN3(\FIFO[3][28] ), .IN4(n6002), 
        .Q(n4463) );
  AO22X1 U4422 ( .IN1(n6763), .IN2(n5998), .IN3(\FIFO[3][29] ), .IN4(n6002), 
        .Q(n4464) );
  AO22X1 U4424 ( .IN1(n6741), .IN2(n5998), .IN3(\FIFO[3][31] ), .IN4(n6002), 
        .Q(n4466) );
  AO21X1 U4425 ( .IN1(n374), .IN2(n263), .IN3(n7361), .Q(n393) );
  AND2X1 U4426 ( .IN1(n394), .IN2(n376), .Q(n263) );
  AO22X1 U4451 ( .IN1(n6818), .IN2(n5991), .IN3(\FIFO[2][24] ), .IN4(n5996), 
        .Q(n4491) );
  AO22X1 U4452 ( .IN1(n6807), .IN2(n5991), .IN3(\FIFO[2][25] ), .IN4(n5996), 
        .Q(n4492) );
  AO22X1 U4453 ( .IN1(n6796), .IN2(n5991), .IN3(\FIFO[2][26] ), .IN4(n5996), 
        .Q(n4493) );
  AO22X1 U4454 ( .IN1(n6785), .IN2(n5991), .IN3(\FIFO[2][27] ), .IN4(n5996), 
        .Q(n4494) );
  AO22X1 U4455 ( .IN1(n6774), .IN2(n5991), .IN3(\FIFO[2][28] ), .IN4(n5996), 
        .Q(n4495) );
  AO22X1 U4456 ( .IN1(n6763), .IN2(n5992), .IN3(\FIFO[2][29] ), .IN4(n5996), 
        .Q(n4496) );
  AO22X1 U4457 ( .IN1(n6752), .IN2(n5991), .IN3(\FIFO[2][30] ), .IN4(n5996), 
        .Q(n4497) );
  AO21X1 U4459 ( .IN1(n374), .IN2(n265), .IN3(n7361), .Q(n395) );
  AND2X1 U4460 ( .IN1(n394), .IN2(n378), .Q(n265) );
  AO22X1 U4461 ( .IN1(n7088), .IN2(n5987), .IN3(\FIFO[1][0] ), .IN4(n5988), 
        .Q(n4499) );
  AO22X1 U4462 ( .IN1(n7071), .IN2(n5987), .IN3(\FIFO[1][1] ), .IN4(n5988), 
        .Q(n4500) );
  AO22X1 U4463 ( .IN1(n7060), .IN2(n5987), .IN3(\FIFO[1][2] ), .IN4(n5988), 
        .Q(n4501) );
  AO22X1 U4464 ( .IN1(n7049), .IN2(n5987), .IN3(\FIFO[1][3] ), .IN4(n5988), 
        .Q(n4502) );
  AO22X1 U4465 ( .IN1(n7038), .IN2(n5987), .IN3(\FIFO[1][4] ), .IN4(n5988), 
        .Q(n4503) );
  AO22X1 U4466 ( .IN1(n7027), .IN2(n5987), .IN3(\FIFO[1][5] ), .IN4(n5988), 
        .Q(n4504) );
  AO22X1 U4468 ( .IN1(n7005), .IN2(n5986), .IN3(\FIFO[1][7] ), .IN4(n5988), 
        .Q(n4506) );
  AO22X1 U4469 ( .IN1(n6994), .IN2(n5986), .IN3(\FIFO[1][8] ), .IN4(n5988), 
        .Q(n4507) );
  AO22X1 U4470 ( .IN1(n6983), .IN2(n5986), .IN3(\FIFO[1][9] ), .IN4(n5988), 
        .Q(n4508) );
  AO22X1 U4471 ( .IN1(n6972), .IN2(n5986), .IN3(\FIFO[1][10] ), .IN4(n5988), 
        .Q(n4509) );
  AO22X1 U4472 ( .IN1(n6961), .IN2(n5986), .IN3(\FIFO[1][11] ), .IN4(n5988), 
        .Q(n4510) );
  AO22X1 U4473 ( .IN1(n6950), .IN2(n5986), .IN3(\FIFO[1][12] ), .IN4(n5989), 
        .Q(n4511) );
  AO22X1 U4474 ( .IN1(n6939), .IN2(n5986), .IN3(\FIFO[1][13] ), .IN4(n5989), 
        .Q(n4512) );
  AO22X1 U4475 ( .IN1(n6928), .IN2(n5985), .IN3(\FIFO[1][14] ), .IN4(n5989), 
        .Q(n4513) );
  AO22X1 U4476 ( .IN1(n6917), .IN2(n5985), .IN3(\FIFO[1][15] ), .IN4(n5989), 
        .Q(n4514) );
  AO22X1 U4477 ( .IN1(n6906), .IN2(n5985), .IN3(\FIFO[1][16] ), .IN4(n5989), 
        .Q(n4515) );
  AO22X1 U4478 ( .IN1(n6895), .IN2(n5985), .IN3(\FIFO[1][17] ), .IN4(n5989), 
        .Q(n4516) );
  AO22X1 U4479 ( .IN1(n6884), .IN2(n5985), .IN3(\FIFO[1][18] ), .IN4(n5989), 
        .Q(n4517) );
  AO22X1 U4480 ( .IN1(n6873), .IN2(n5985), .IN3(\FIFO[1][19] ), .IN4(n5989), 
        .Q(n4518) );
  AO22X1 U4481 ( .IN1(n6862), .IN2(n5985), .IN3(\FIFO[1][20] ), .IN4(n5989), 
        .Q(n4519) );
  AO22X1 U4482 ( .IN1(n6851), .IN2(n5987), .IN3(\FIFO[1][21] ), .IN4(n5989), 
        .Q(n4520) );
  AO22X1 U4484 ( .IN1(n6829), .IN2(n5985), .IN3(\FIFO[1][23] ), .IN4(n5989), 
        .Q(n4522) );
  AO22X1 U4485 ( .IN1(n6818), .IN2(n396), .IN3(\FIFO[1][24] ), .IN4(n5990), 
        .Q(n4523) );
  AO22X1 U4486 ( .IN1(n6807), .IN2(n396), .IN3(\FIFO[1][25] ), .IN4(n5990), 
        .Q(n4524) );
  AO22X1 U4487 ( .IN1(n6796), .IN2(n396), .IN3(\FIFO[1][26] ), .IN4(n5990), 
        .Q(n4525) );
  AO22X1 U4488 ( .IN1(n6785), .IN2(n5987), .IN3(\FIFO[1][27] ), .IN4(n5990), 
        .Q(n4526) );
  AO22X1 U4489 ( .IN1(n6774), .IN2(n5986), .IN3(\FIFO[1][28] ), .IN4(n5990), 
        .Q(n4527) );
  AO22X1 U4490 ( .IN1(n6763), .IN2(n5987), .IN3(\FIFO[1][29] ), .IN4(n5990), 
        .Q(n4528) );
  AO22X1 U4491 ( .IN1(n6752), .IN2(n5986), .IN3(\FIFO[1][30] ), .IN4(n5990), 
        .Q(n4529) );
  AO22X1 U4492 ( .IN1(n6741), .IN2(n5985), .IN3(\FIFO[1][31] ), .IN4(n5990), 
        .Q(n4530) );
  AO21X1 U4493 ( .IN1(n374), .IN2(n267), .IN3(n7361), .Q(n396) );
  AND2X1 U4494 ( .IN1(n394), .IN2(n380), .Q(n267) );
  AO22X1 U4495 ( .IN1(n7088), .IN2(n5980), .IN3(n5982), .IN4(\FIFO[0][0] ), 
        .Q(n4531) );
  AO22X1 U4497 ( .IN1(n7071), .IN2(n5979), .IN3(n5982), .IN4(\FIFO[0][1] ), 
        .Q(n4532) );
  AO22X1 U4499 ( .IN1(n7060), .IN2(n5981), .IN3(n5982), .IN4(\FIFO[0][2] ), 
        .Q(n4533) );
  AO22X1 U4501 ( .IN1(n7049), .IN2(n5980), .IN3(n5982), .IN4(\FIFO[0][3] ), 
        .Q(n4534) );
  AO22X1 U4503 ( .IN1(n7038), .IN2(n5979), .IN3(n5982), .IN4(\FIFO[0][4] ), 
        .Q(n4535) );
  AO22X1 U4505 ( .IN1(n7027), .IN2(n5981), .IN3(n5982), .IN4(\FIFO[0][5] ), 
        .Q(n4536) );
  AO22X1 U4507 ( .IN1(n7016), .IN2(n5980), .IN3(n5982), .IN4(\FIFO[0][6] ), 
        .Q(n4537) );
  AO22X1 U4509 ( .IN1(n7005), .IN2(n5980), .IN3(n5982), .IN4(\FIFO[0][7] ), 
        .Q(n4538) );
  AO22X1 U4511 ( .IN1(n6994), .IN2(n5979), .IN3(n5982), .IN4(\FIFO[0][8] ), 
        .Q(n4539) );
  AO22X1 U4513 ( .IN1(n6983), .IN2(n5981), .IN3(n5982), .IN4(\FIFO[0][9] ), 
        .Q(n4540) );
  AO22X1 U4515 ( .IN1(n6972), .IN2(n5980), .IN3(n5982), .IN4(\FIFO[0][10] ), 
        .Q(n4541) );
  AO22X1 U4519 ( .IN1(n6950), .IN2(n5980), .IN3(n5983), .IN4(\FIFO[0][12] ), 
        .Q(n4543) );
  AO22X1 U4521 ( .IN1(n6939), .IN2(n5979), .IN3(n5983), .IN4(\FIFO[0][13] ), 
        .Q(n4544) );
  AO22X1 U4523 ( .IN1(n6928), .IN2(n5979), .IN3(n5983), .IN4(\FIFO[0][14] ), 
        .Q(n4545) );
  AO22X1 U4525 ( .IN1(n6917), .IN2(n5981), .IN3(n5983), .IN4(\FIFO[0][15] ), 
        .Q(n4546) );
  AO22X1 U4527 ( .IN1(n6906), .IN2(n5980), .IN3(n5983), .IN4(\FIFO[0][16] ), 
        .Q(n4547) );
  AO22X1 U4529 ( .IN1(n6895), .IN2(n5979), .IN3(n5983), .IN4(\FIFO[0][17] ), 
        .Q(n4548) );
  AO22X1 U4531 ( .IN1(n6884), .IN2(n5981), .IN3(n5983), .IN4(\FIFO[0][18] ), 
        .Q(n4549) );
  AO22X1 U4533 ( .IN1(n6873), .IN2(n5980), .IN3(n5983), .IN4(\FIFO[0][19] ), 
        .Q(n4550) );
  AO22X1 U4535 ( .IN1(n6862), .IN2(n5979), .IN3(n5983), .IN4(\FIFO[0][20] ), 
        .Q(n4551) );
  AO22X1 U4537 ( .IN1(n6851), .IN2(n5981), .IN3(n5983), .IN4(\FIFO[0][21] ), 
        .Q(n4552) );
  AO22X1 U4539 ( .IN1(n6840), .IN2(n5981), .IN3(n5983), .IN4(\FIFO[0][22] ), 
        .Q(n4553) );
  AO22X1 U4543 ( .IN1(n6818), .IN2(n397), .IN3(n5984), .IN4(\FIFO[0][24] ), 
        .Q(n4555) );
  AO22X1 U4545 ( .IN1(n6807), .IN2(n397), .IN3(n5984), .IN4(\FIFO[0][25] ), 
        .Q(n4556) );
  AO22X1 U4547 ( .IN1(n6796), .IN2(n397), .IN3(n5984), .IN4(\FIFO[0][26] ), 
        .Q(n4557) );
  AO22X1 U4549 ( .IN1(n6785), .IN2(n5979), .IN3(n5984), .IN4(\FIFO[0][27] ), 
        .Q(n4558) );
  AO22X1 U4551 ( .IN1(n6774), .IN2(n5979), .IN3(n5984), .IN4(\FIFO[0][28] ), 
        .Q(n4559) );
  AO22X1 U4553 ( .IN1(n6763), .IN2(n5981), .IN3(n5984), .IN4(\FIFO[0][29] ), 
        .Q(n4560) );
  AO22X1 U4555 ( .IN1(n6752), .IN2(n5981), .IN3(n5984), .IN4(\FIFO[0][30] ), 
        .Q(n4561) );
  AO22X1 U4557 ( .IN1(n6741), .IN2(n5980), .IN3(n5984), .IN4(\FIFO[0][31] ), 
        .Q(n4562) );
  AO21X1 U4558 ( .IN1(n374), .IN2(n269), .IN3(n7361), .Q(n397) );
  AND2X1 U4559 ( .IN1(n394), .IN2(n382), .Q(n269) );
  AO22X1 U4565 ( .IN1(\FIFO[0][27] ), .IN2(n7103), .IN3(N223), .IN4(n204), .Q(
        N280) );
  AO22X1 U4566 ( .IN1(\FIFO[0][26] ), .IN2(n7101), .IN3(N224), .IN4(n204), .Q(
        N279) );
  AO22X1 U4567 ( .IN1(\FIFO[0][25] ), .IN2(n7102), .IN3(N225), .IN4(n204), .Q(
        N278) );
  AO22X1 U4568 ( .IN1(\FIFO[0][24] ), .IN2(n7103), .IN3(N226), .IN4(n204), .Q(
        N277) );
  AO22X1 U4569 ( .IN1(\FIFO[0][23] ), .IN2(n7101), .IN3(N227), .IN4(n7100), 
        .Q(N276) );
  AO22X1 U4570 ( .IN1(\FIFO[0][22] ), .IN2(n7102), .IN3(N228), .IN4(n7100), 
        .Q(N275) );
  AO22X1 U4571 ( .IN1(\FIFO[0][21] ), .IN2(n7103), .IN3(N229), .IN4(n7100), 
        .Q(N274) );
  AO22X1 U4572 ( .IN1(\FIFO[0][20] ), .IN2(n7101), .IN3(N230), .IN4(n7100), 
        .Q(N273) );
  AO22X1 U4573 ( .IN1(\FIFO[0][19] ), .IN2(n7101), .IN3(N231), .IN4(n7100), 
        .Q(N272) );
  AO22X1 U4574 ( .IN1(\FIFO[0][18] ), .IN2(n7101), .IN3(N232), .IN4(n7100), 
        .Q(N271) );
  AO22X1 U4575 ( .IN1(\FIFO[0][17] ), .IN2(n7101), .IN3(N233), .IN4(n7100), 
        .Q(N270) );
  AO22X1 U4576 ( .IN1(\FIFO[0][16] ), .IN2(n7101), .IN3(N234), .IN4(n7100), 
        .Q(N269) );
  AO22X1 U4577 ( .IN1(\FIFO[0][15] ), .IN2(n7101), .IN3(N235), .IN4(n7100), 
        .Q(N268) );
  AO22X1 U4578 ( .IN1(\FIFO[0][14] ), .IN2(n7101), .IN3(N236), .IN4(n7100), 
        .Q(N267) );
  AO22X1 U4579 ( .IN1(\FIFO[0][13] ), .IN2(n7102), .IN3(N237), .IN4(n7100), 
        .Q(N266) );
  AO22X1 U4580 ( .IN1(\FIFO[0][12] ), .IN2(n7102), .IN3(N238), .IN4(n7100), 
        .Q(N265) );
  AO22X1 U4581 ( .IN1(\FIFO[0][11] ), .IN2(n7102), .IN3(N239), .IN4(n7099), 
        .Q(N264) );
  AO22X1 U4582 ( .IN1(\FIFO[0][10] ), .IN2(n7102), .IN3(N240), .IN4(n7099), 
        .Q(N263) );
  AO22X1 U4583 ( .IN1(\FIFO[0][9] ), .IN2(n7102), .IN3(N241), .IN4(n7099), .Q(
        N262) );
  AO22X1 U4584 ( .IN1(\FIFO[0][8] ), .IN2(n7102), .IN3(N242), .IN4(n7099), .Q(
        N261) );
  AO22X1 U4585 ( .IN1(\FIFO[0][7] ), .IN2(n7102), .IN3(N243), .IN4(n7099), .Q(
        N260) );
  AO22X1 U4586 ( .IN1(\FIFO[0][6] ), .IN2(n7103), .IN3(N244), .IN4(n7099), .Q(
        N259) );
  AO22X1 U4587 ( .IN1(\FIFO[0][5] ), .IN2(n7103), .IN3(N245), .IN4(n7099), .Q(
        N258) );
  AO22X1 U4588 ( .IN1(\FIFO[0][4] ), .IN2(n7103), .IN3(N246), .IN4(n7099), .Q(
        N257) );
  AO22X1 U4589 ( .IN1(\FIFO[0][3] ), .IN2(n7103), .IN3(N247), .IN4(n7099), .Q(
        N256) );
  AO22X1 U4590 ( .IN1(\FIFO[0][2] ), .IN2(n7103), .IN3(N248), .IN4(n7099), .Q(
        N255) );
  AO22X1 U4591 ( .IN1(\FIFO[0][1] ), .IN2(n7103), .IN3(N249), .IN4(n7099), .Q(
        N254) );
  AO22X1 U4592 ( .IN1(\FIFO[0][0] ), .IN2(n7103), .IN3(N250), .IN4(n7099), .Q(
        N253) );
  OR3X1 U4594 ( .IN1(rden), .IN2(rdaddr[7]), .IN3(N21), .Q(n401) );
  OR4X1 U4595 ( .IN1(N15), .IN2(N16), .IN3(N17), .IN4(N18), .Q(n400) );
  AND2X4 U3 ( .IN1(n374), .IN2(n259), .Q(n1) );
  OR2X4 U4 ( .IN1(n1), .IN2(n7361), .Q(n391) );
  AND2X4 U5 ( .IN1(n389), .IN2(n380), .Q(n259) );
  DELLN1X2 U6 ( .INP(n391), .Z(n6009) );
  DELLN1X2 U7 ( .INP(n391), .Z(n6010) );
  DELLN1X2 U8 ( .INP(n391), .Z(n6011) );
  MUX21X1 U9 ( .IN1(\FIFO[5][20] ), .IN2(n51), .S(n391), .Q(n4391) );
  MUX21X1 U10 ( .IN1(\FIFO[5][9] ), .IN2(n27), .S(n391), .Q(n4380) );
  AND2X4 U11 ( .IN1(n374), .IN2(n257), .Q(n2) );
  OR2X4 U12 ( .IN1(n2), .IN2(n7361), .Q(n390) );
  AND2X4 U13 ( .IN1(n389), .IN2(n378), .Q(n257) );
  DELLN1X2 U14 ( .INP(n390), .Z(n6015) );
  DELLN1X2 U15 ( .INP(n390), .Z(n6016) );
  DELLN1X2 U16 ( .INP(n390), .Z(n6017) );
  MUX21X1 U17 ( .IN1(\FIFO[6][19] ), .IN2(n23), .S(n390), .Q(n4358) );
  MUX21X1 U18 ( .IN1(\FIFO[6][8] ), .IN2(n50), .S(n390), .Q(n4347) );
  AND2X4 U19 ( .IN1(n374), .IN2(n251), .Q(n3) );
  OR2X4 U20 ( .IN1(n3), .IN2(n7361), .Q(n386) );
  AND2X4 U21 ( .IN1(n384), .IN2(n380), .Q(n251) );
  DELLN1X2 U22 ( .INP(n386), .Z(n6033) );
  DELLN1X2 U23 ( .INP(n386), .Z(n6034) );
  DELLN1X2 U24 ( .INP(n386), .Z(n6035) );
  MUX21X1 U25 ( .IN1(\FIFO[9][18] ), .IN2(n24), .S(n386), .Q(n4261) );
  MUX21X1 U26 ( .IN1(\FIFO[9][7] ), .IN2(n42), .S(n386), .Q(n4250) );
  AND2X4 U27 ( .IN1(n374), .IN2(n249), .Q(n4) );
  OR2X4 U28 ( .IN1(n4), .IN2(n7361), .Q(n385) );
  AND2X4 U29 ( .IN1(n384), .IN2(n378), .Q(n249) );
  DELLN1X2 U30 ( .INP(n385), .Z(n6039) );
  DELLN1X2 U31 ( .INP(n385), .Z(n6040) );
  DELLN1X2 U32 ( .INP(n385), .Z(n6041) );
  MUX21X1 U33 ( .IN1(\FIFO[10][17] ), .IN2(n28), .S(n385), .Q(n4228) );
  MUX21X1 U34 ( .IN1(\FIFO[10][5] ), .IN2(n44), .S(n385), .Q(n4216) );
  AND2X4 U35 ( .IN1(n374), .IN2(n247), .Q(n5) );
  OR2X4 U36 ( .IN1(n5), .IN2(n7361), .Q(n383) );
  AND2X4 U37 ( .IN1(n384), .IN2(n376), .Q(n247) );
  DELLN1X2 U38 ( .INP(n383), .Z(n6045) );
  DELLN1X2 U39 ( .INP(n383), .Z(n6046) );
  DELLN1X2 U40 ( .INP(n383), .Z(n6047) );
  MUX21X1 U41 ( .IN1(\FIFO[11][16] ), .IN2(n29), .S(n383), .Q(n4195) );
  MUX21X1 U42 ( .IN1(\FIFO[11][4] ), .IN2(n45), .S(n383), .Q(n4183) );
  AND2X4 U43 ( .IN1(n374), .IN2(n241), .Q(n6) );
  OR2X4 U44 ( .IN1(n6), .IN2(n7361), .Q(n377) );
  AND2X4 U45 ( .IN1(n378), .IN2(n375), .Q(n241) );
  DELLN1X2 U46 ( .INP(n377), .Z(n6063) );
  DELLN1X2 U47 ( .INP(n377), .Z(n6064) );
  DELLN1X2 U48 ( .INP(n377), .Z(n6065) );
  MUX21X1 U49 ( .IN1(\FIFO[14][15] ), .IN2(n30), .S(n377), .Q(n4098) );
  MUX21X1 U50 ( .IN1(\FIFO[14][3] ), .IN2(n46), .S(n377), .Q(n4086) );
  AND2X4 U51 ( .IN1(n374), .IN2(n238), .Q(n7) );
  OR2X4 U52 ( .IN1(n7), .IN2(n7361), .Q(n373) );
  AND2X4 U53 ( .IN1(n375), .IN2(n376), .Q(n238) );
  DELLN1X2 U54 ( .INP(n373), .Z(n6069) );
  DELLN1X2 U55 ( .INP(n373), .Z(n6070) );
  DELLN1X2 U56 ( .INP(n373), .Z(n6071) );
  MUX21X1 U57 ( .IN1(\FIFO[15][14] ), .IN2(n31), .S(n373), .Q(n4065) );
  MUX21X1 U58 ( .IN1(\FIFO[15][2] ), .IN2(n47), .S(n373), .Q(n4053) );
  OR2X4 U59 ( .IN1(wren), .IN2(n5973), .Q(n8) );
  MUX21X1 U60 ( .IN1(\FIFO[0][28] ), .IN2(N222), .S(n204), .Q(N281) );
  MUX21X1 U61 ( .IN1(\FIFO[0][29] ), .IN2(N221), .S(n204), .Q(N282) );
  MUX21X1 U62 ( .IN1(\FIFO[0][30] ), .IN2(N220), .S(n204), .Q(N283) );
  MUX21X1 U63 ( .IN1(\FIFO[0][31] ), .IN2(N219), .S(n204), .Q(n464) );
  MUX21X1 U64 ( .IN1(\FIFO[115][6] ), .IN2(n43), .S(n262), .Q(n857) );
  MUX21X1 U65 ( .IN1(\FIFO[113][7] ), .IN2(n42), .S(n266), .Q(n922) );
  MUX21X1 U66 ( .IN1(\FIFO[108][8] ), .IN2(n50), .S(n275), .Q(n1083) );
  MUX21X1 U67 ( .IN1(\FIFO[103][12] ), .IN2(n33), .S(n280), .Q(n1247) );
  MUX21X1 U68 ( .IN1(\FIFO[102][1] ), .IN2(n48), .S(n281), .Q(n1268) );
  MUX21X1 U69 ( .IN1(\FIFO[98][13] ), .IN2(n32), .S(n285), .Q(n1408) );
  MUX21X1 U70 ( .IN1(\FIFO[97][0] ), .IN2(n49), .S(n286), .Q(n1427) );
  MUX21X1 U71 ( .IN1(\FIFO[97][14] ), .IN2(n31), .S(n286), .Q(n1441) );
  MUX21X1 U72 ( .IN1(\FIFO[94][1] ), .IN2(n48), .S(n290), .Q(n1524) );
  MUX21X1 U73 ( .IN1(\FIFO[94][15] ), .IN2(n30), .S(n290), .Q(n1538) );
  MUX21X1 U74 ( .IN1(\FIFO[93][2] ), .IN2(n47), .S(n291), .Q(n1557) );
  MUX21X1 U75 ( .IN1(\FIFO[93][17] ), .IN2(n28), .S(n291), .Q(n1572) );
  MUX21X1 U76 ( .IN1(\FIFO[89][3] ), .IN2(n46), .S(n295), .Q(n1686) );
  MUX21X1 U77 ( .IN1(\FIFO[89][16] ), .IN2(n29), .S(n295), .Q(n1699) );
  MUX21X1 U78 ( .IN1(\FIFO[88][4] ), .IN2(n45), .S(n296), .Q(n1719) );
  MUX21X1 U79 ( .IN1(\FIFO[84][5] ), .IN2(n44), .S(n300), .Q(n1848) );
  MUX21X1 U80 ( .IN1(\FIFO[84][18] ), .IN2(n24), .S(n300), .Q(n1861) );
  MUX21X1 U81 ( .IN1(\FIFO[83][6] ), .IN2(n43), .S(n301), .Q(n1881) );
  MUX21X1 U82 ( .IN1(\FIFO[83][20] ), .IN2(n51), .S(n301), .Q(n1895) );
  MUX21X1 U83 ( .IN1(\FIFO[77][7] ), .IN2(n42), .S(n308), .Q(n2074) );
  MUX21X1 U84 ( .IN1(\FIFO[77][19] ), .IN2(n23), .S(n308), .Q(n2086) );
  MUX21X1 U85 ( .IN1(\FIFO[76][8] ), .IN2(n50), .S(n309), .Q(n2107) );
  MUX21X1 U86 ( .IN1(\FIFO[76][21] ), .IN2(n22), .S(n309), .Q(n2120) );
  MUX21X1 U87 ( .IN1(\FIFO[72][9] ), .IN2(n27), .S(n313), .Q(n2236) );
  MUX21X1 U88 ( .IN1(\FIFO[72][22] ), .IN2(n21), .S(n313), .Q(n2249) );
  MUX21X1 U89 ( .IN1(\FIFO[71][10] ), .IN2(n26), .S(n314), .Q(n2269) );
  MUX21X1 U90 ( .IN1(\FIFO[71][23] ), .IN2(n20), .S(n314), .Q(n2282) );
  MUX21X1 U91 ( .IN1(\FIFO[67][12] ), .IN2(n33), .S(n318), .Q(n2399) );
  MUX21X1 U92 ( .IN1(\FIFO[66][4] ), .IN2(n45), .S(n319), .Q(n2423) );
  MUX21X1 U93 ( .IN1(\FIFO[66][13] ), .IN2(n32), .S(n319), .Q(n2432) );
  MUX21X1 U94 ( .IN1(\FIFO[63][9] ), .IN2(n27), .S(n322), .Q(n2524) );
  MUX21X1 U95 ( .IN1(\FIFO[63][14] ), .IN2(n31), .S(n322), .Q(n2529) );
  MUX21X1 U96 ( .IN1(\FIFO[62][15] ), .IN2(n30), .S(n324), .Q(n2562) );
  MUX21X1 U97 ( .IN1(\FIFO[58][10] ), .IN2(n26), .S(n328), .Q(n2685) );
  MUX21X1 U98 ( .IN1(\FIFO[58][16] ), .IN2(n29), .S(n328), .Q(n2691) );
  MUX21X1 U99 ( .IN1(\FIFO[57][2] ), .IN2(n47), .S(n329), .Q(n2709) );
  MUX21X1 U100 ( .IN1(\FIFO[57][17] ), .IN2(n28), .S(n329), .Q(n2724) );
  MUX21X1 U101 ( .IN1(\FIFO[53][18] ), .IN2(n24), .S(n333), .Q(n2853) );
  MUX21X1 U102 ( .IN1(\FIFO[52][5] ), .IN2(n44), .S(n334), .Q(n2872) );
  MUX21X1 U103 ( .IN1(\FIFO[52][19] ), .IN2(n23), .S(n334), .Q(n2886) );
  MUX21X1 U104 ( .IN1(\FIFO[48][11] ), .IN2(n25), .S(n338), .Q(n3006) );
  MUX21X1 U105 ( .IN1(\FIFO[48][20] ), .IN2(n51), .S(n338), .Q(n3015) );
  MUX21X1 U106 ( .IN1(\FIFO[44][0] ), .IN2(n49), .S(n343), .Q(n3123) );
  MUX21X1 U107 ( .IN1(\FIFO[44][21] ), .IN2(n22), .S(n343), .Q(n3144) );
  MUX21X1 U108 ( .IN1(\FIFO[43][1] ), .IN2(n48), .S(n344), .Q(n3156) );
  MUX21X1 U109 ( .IN1(\FIFO[43][22] ), .IN2(n21), .S(n344), .Q(n3177) );
  MUX21X1 U110 ( .IN1(\FIFO[42][4] ), .IN2(n45), .S(n345), .Q(n3191) );
  MUX21X1 U111 ( .IN1(\FIFO[41][8] ), .IN2(n50), .S(n346), .Q(n3227) );
  MUX21X1 U112 ( .IN1(\FIFO[40][9] ), .IN2(n27), .S(n347), .Q(n3260) );
  MUX21X1 U113 ( .IN1(\FIFO[39][14] ), .IN2(n31), .S(n348), .Q(n3297) );
  MUX21X1 U114 ( .IN1(\FIFO[39][23] ), .IN2(n20), .S(n348), .Q(n3306) );
  MUX21X1 U115 ( .IN1(\FIFO[38][16] ), .IN2(n29), .S(n349), .Q(n3331) );
  MUX21X1 U116 ( .IN1(\FIFO[38][24] ), .IN2(n41), .S(n349), .Q(n3339) );
  MUX21X1 U117 ( .IN1(\FIFO[37][10] ), .IN2(n26), .S(n350), .Q(n3357) );
  MUX21X1 U118 ( .IN1(\FIFO[36][12] ), .IN2(n33), .S(n351), .Q(n3391) );
  MUX21X1 U119 ( .IN1(\FIFO[35][14] ), .IN2(n31), .S(n352), .Q(n3425) );
  MUX21X1 U120 ( .IN1(\FIFO[34][11] ), .IN2(n25), .S(n353), .Q(n3454) );
  MUX21X1 U121 ( .IN1(\FIFO[34][17] ), .IN2(n28), .S(n353), .Q(n3460) );
  MUX21X1 U122 ( .IN1(\FIFO[34][25] ), .IN2(n40), .S(n353), .Q(n3468) );
  MUX21X1 U123 ( .IN1(\FIFO[33][18] ), .IN2(n24), .S(n354), .Q(n3493) );
  MUX21X1 U124 ( .IN1(\FIFO[33][26] ), .IN2(n39), .S(n354), .Q(n3501) );
  MUX21X1 U125 ( .IN1(\FIFO[32][15] ), .IN2(n30), .S(n355), .Q(n3522) );
  MUX21X1 U126 ( .IN1(\FIFO[31][0] ), .IN2(n49), .S(n356), .Q(n3539) );
  MUX21X1 U127 ( .IN1(\FIFO[31][19] ), .IN2(n23), .S(n356), .Q(n3558) );
  MUX21X1 U128 ( .IN1(\FIFO[31][27] ), .IN2(n38), .S(n356), .Q(n3566) );
  MUX21X1 U129 ( .IN1(\FIFO[30][1] ), .IN2(n48), .S(n358), .Q(n3572) );
  MUX21X1 U130 ( .IN1(\FIFO[29][2] ), .IN2(n47), .S(n359), .Q(n3605) );
  MUX21X1 U131 ( .IN1(\FIFO[27][4] ), .IN2(n45), .S(n361), .Q(n3671) );
  MUX21X1 U132 ( .IN1(\FIFO[27][20] ), .IN2(n51), .S(n361), .Q(n3687) );
  MUX21X1 U133 ( .IN1(\FIFO[27][28] ), .IN2(n37), .S(n361), .Q(n3695) );
  MUX21X1 U134 ( .IN1(\FIFO[26][5] ), .IN2(n44), .S(n362), .Q(n3704) );
  MUX21X1 U135 ( .IN1(\FIFO[26][21] ), .IN2(n22), .S(n362), .Q(n3720) );
  MUX21X1 U136 ( .IN1(\FIFO[26][29] ), .IN2(n36), .S(n362), .Q(n3728) );
  MUX21X1 U137 ( .IN1(\FIFO[24][7] ), .IN2(n42), .S(n364), .Q(n3770) );
  MUX21X1 U138 ( .IN1(\FIFO[23][8] ), .IN2(n50), .S(n365), .Q(n3803) );
  MUX21X1 U139 ( .IN1(\FIFO[22][9] ), .IN2(n27), .S(n366), .Q(n3836) );
  MUX21X1 U140 ( .IN1(\FIFO[22][22] ), .IN2(n21), .S(n366), .Q(n3849) );
  MUX21X1 U141 ( .IN1(\FIFO[22][30] ), .IN2(n35), .S(n366), .Q(n3857) );
  MUX21X1 U142 ( .IN1(\FIFO[21][10] ), .IN2(n26), .S(n367), .Q(n3869) );
  MUX21X1 U143 ( .IN1(\FIFO[21][23] ), .IN2(n20), .S(n367), .Q(n3882) );
  MUX21X1 U144 ( .IN1(\FIFO[21][31] ), .IN2(n34), .S(n367), .Q(n3890) );
  MUX21X1 U145 ( .IN1(\FIFO[20][11] ), .IN2(n25), .S(n368), .Q(n3902) );
  MUX21X1 U146 ( .IN1(\FIFO[17][11] ), .IN2(n25), .S(n371), .Q(n3998) );
  MUX21X1 U147 ( .IN1(\FIFO[17][16] ), .IN2(n29), .S(n371), .Q(n4003) );
  MUX21X1 U148 ( .IN1(\FIFO[17][24] ), .IN2(n41), .S(n371), .Q(n4011) );
  MUX21X1 U149 ( .IN1(\FIFO[16][5] ), .IN2(n44), .S(n372), .Q(n4024) );
  MUX21X1 U150 ( .IN1(\FIFO[16][17] ), .IN2(n28), .S(n372), .Q(n4036) );
  MUX21X1 U151 ( .IN1(\FIFO[16][25] ), .IN2(n40), .S(n372), .Q(n4044) );
  MUX21X1 U152 ( .IN1(\FIFO[13][6] ), .IN2(n43), .S(n379), .Q(n4121) );
  MUX21X1 U153 ( .IN1(\FIFO[13][18] ), .IN2(n24), .S(n379), .Q(n4133) );
  MUX21X1 U154 ( .IN1(\FIFO[13][26] ), .IN2(n39), .S(n379), .Q(n4141) );
  MUX21X1 U155 ( .IN1(\FIFO[12][7] ), .IN2(n42), .S(n381), .Q(n4154) );
  MUX21X1 U156 ( .IN1(\FIFO[12][19] ), .IN2(n23), .S(n381), .Q(n4166) );
  MUX21X1 U157 ( .IN1(\FIFO[12][27] ), .IN2(n38), .S(n381), .Q(n4174) );
  MUX21X1 U158 ( .IN1(\FIFO[8][13] ), .IN2(n32), .S(n387), .Q(n4288) );
  MUX21X1 U159 ( .IN1(\FIFO[8][20] ), .IN2(n51), .S(n387), .Q(n4295) );
  MUX21X1 U160 ( .IN1(\FIFO[8][28] ), .IN2(n37), .S(n387), .Q(n4303) );
  MUX21X1 U161 ( .IN1(\FIFO[7][2] ), .IN2(n47), .S(n388), .Q(n4309) );
  MUX21X1 U162 ( .IN1(\FIFO[7][21] ), .IN2(n22), .S(n388), .Q(n4328) );
  MUX21X1 U163 ( .IN1(\FIFO[7][29] ), .IN2(n36), .S(n388), .Q(n4336) );
  MUX21X1 U164 ( .IN1(\FIFO[3][15] ), .IN2(n30), .S(n393), .Q(n4450) );
  MUX21X1 U165 ( .IN1(\FIFO[3][22] ), .IN2(n21), .S(n393), .Q(n4457) );
  MUX21X1 U166 ( .IN1(\FIFO[3][30] ), .IN2(n35), .S(n393), .Q(n4465) );
  MUX21X1 U167 ( .IN1(\FIFO[2][3] ), .IN2(n46), .S(n395), .Q(n4470) );
  MUX21X1 U168 ( .IN1(\FIFO[2][23] ), .IN2(n20), .S(n395), .Q(n4490) );
  MUX21X1 U169 ( .IN1(\FIFO[2][31] ), .IN2(n34), .S(n395), .Q(n4498) );
  NAND2X1 U170 ( .IN1(n11), .IN2(n7356), .QN(n63) );
  NAND2X1 U171 ( .IN1(n9), .IN2(n7340), .QN(n74) );
  NAND2X1 U172 ( .IN1(n10), .IN2(n7348), .QN(n81) );
  NAND2X1 U173 ( .IN1(n15), .IN2(n7358), .QN(n84) );
  NAND2X1 U174 ( .IN1(n14), .IN2(n7355), .QN(n64) );
  NAND2X1 U175 ( .IN1(n18), .IN2(n7344), .QN(n76) );
  NAND2X1 U176 ( .IN1(n12), .IN2(n7340), .QN(n75) );
  NAND2X1 U177 ( .IN1(n16), .IN2(n7351), .QN(n77) );
  NAND2X1 U178 ( .IN1(n13), .IN2(n7348), .QN(n83) );
  NAND2X1 U179 ( .IN1(n7355), .IN2(\FIFO[0][3] ), .QN(n89) );
  NAND2X1 U180 ( .IN1(n7357), .IN2(\FIFO[0][18] ), .QN(n104) );
  NAND2X1 U181 ( .IN1(n7356), .IN2(\FIFO[0][21] ), .QN(n107) );
  NAND2X1 U182 ( .IN1(n19), .IN2(n7354), .QN(n85) );
  MUX21X2 U183 ( .IN1(\FIFO[28][12] ), .IN2(n33), .S(n360), .Q(n3647) );
  MUX21X2 U184 ( .IN1(\FIFO[25][13] ), .IN2(n32), .S(n363), .Q(n3744) );
  MUX21X2 U185 ( .IN1(\FIFO[19][0] ), .IN2(n49), .S(n369), .Q(n3923) );
  MUX21X2 U186 ( .IN1(\FIFO[18][1] ), .IN2(n48), .S(n370), .Q(n3956) );
  MUX21X2 U187 ( .IN1(\FIFO[4][10] ), .IN2(n26), .S(n392), .Q(n4413) );
  MUX21X2 U188 ( .IN1(\FIFO[1][6] ), .IN2(n43), .S(n396), .Q(n4505) );
  MUX21X2 U189 ( .IN1(\FIFO[0][11] ), .IN2(n25), .S(n397), .Q(n4542) );
  AO21X1 U190 ( .IN1(n323), .IN2(n243), .IN3(n7359), .Q(n325) );
  NAND2X1 U191 ( .IN1(n7355), .IN2(\FIFO[0][4] ), .QN(n90) );
  NAND2X1 U192 ( .IN1(n7354), .IN2(\FIFO[0][5] ), .QN(n91) );
  NAND2X1 U193 ( .IN1(n17), .IN2(n7339), .QN(n65) );
  NAND2X1 U194 ( .IN1(n7357), .IN2(\FIFO[0][19] ), .QN(n105) );
  NAND2X1 U195 ( .IN1(n7353), .IN2(\FIFO[0][26] ), .QN(n112) );
  NAND2X1 U196 ( .IN1(n7356), .IN2(\FIFO[0][28] ), .QN(n114) );
  MUX21X2 U197 ( .IN1(\FIFO[28][3] ), .IN2(n46), .S(n360), .Q(n3638) );
  MUX21X2 U198 ( .IN1(\FIFO[25][6] ), .IN2(n43), .S(n363), .Q(n3737) );
  MUX21X2 U199 ( .IN1(\FIFO[19][12] ), .IN2(n33), .S(n369), .Q(n3935) );
  MUX21X2 U200 ( .IN1(\FIFO[18][13] ), .IN2(n32), .S(n370), .Q(n3968) );
  MUX21X2 U201 ( .IN1(\FIFO[4][21] ), .IN2(n22), .S(n392), .Q(n4424) );
  MUX21X2 U202 ( .IN1(\FIFO[1][22] ), .IN2(n21), .S(n396), .Q(n4521) );
  MUX21X2 U203 ( .IN1(\FIFO[0][23] ), .IN2(n20), .S(n397), .Q(n4554) );
  AND2X4 U204 ( .IN1(dataIn[23]), .IN2(n5978), .Q(n20) );
  AND2X4 U205 ( .IN1(dataIn[22]), .IN2(n5976), .Q(n21) );
  AND2X4 U206 ( .IN1(dataIn[21]), .IN2(n5978), .Q(n22) );
  AND2X4 U207 ( .IN1(dataIn[19]), .IN2(n5976), .Q(n23) );
  AND2X4 U208 ( .IN1(dataIn[18]), .IN2(n5977), .Q(n24) );
  AND2X4 U209 ( .IN1(dataIn[11]), .IN2(n5976), .Q(n25) );
  AND2X4 U210 ( .IN1(dataIn[10]), .IN2(n5977), .Q(n26) );
  AND2X4 U211 ( .IN1(dataIn[9]), .IN2(n5978), .Q(n27) );
  AND2X4 U212 ( .IN1(dataIn[17]), .IN2(n5976), .Q(n28) );
  AND2X4 U213 ( .IN1(dataIn[16]), .IN2(n5977), .Q(n29) );
  AND2X4 U214 ( .IN1(dataIn[15]), .IN2(n5978), .Q(n30) );
  AND2X4 U215 ( .IN1(dataIn[14]), .IN2(n5976), .Q(n31) );
  AND2X4 U216 ( .IN1(dataIn[13]), .IN2(n5978), .Q(n32) );
  AND2X4 U217 ( .IN1(dataIn[12]), .IN2(n5976), .Q(n33) );
  AND2X4 U218 ( .IN1(dataIn[31]), .IN2(n5976), .Q(n34) );
  AND2X4 U219 ( .IN1(dataIn[30]), .IN2(n5977), .Q(n35) );
  AND2X4 U220 ( .IN1(dataIn[29]), .IN2(n5978), .Q(n36) );
  AND2X4 U221 ( .IN1(dataIn[28]), .IN2(n5976), .Q(n37) );
  AND2X4 U222 ( .IN1(dataIn[27]), .IN2(n5977), .Q(n38) );
  AND2X4 U223 ( .IN1(dataIn[26]), .IN2(n5976), .Q(n39) );
  AND2X4 U224 ( .IN1(dataIn[25]), .IN2(n5977), .Q(n40) );
  AND2X4 U225 ( .IN1(dataIn[24]), .IN2(n5978), .Q(n41) );
  AND2X4 U226 ( .IN1(dataIn[7]), .IN2(n5977), .Q(n42) );
  AND2X4 U227 ( .IN1(dataIn[6]), .IN2(n5976), .Q(n43) );
  AND2X4 U228 ( .IN1(dataIn[5]), .IN2(n5978), .Q(n44) );
  AND2X4 U229 ( .IN1(dataIn[4]), .IN2(n5976), .Q(n45) );
  AND2X4 U230 ( .IN1(dataIn[3]), .IN2(n5978), .Q(n46) );
  AND2X4 U231 ( .IN1(dataIn[2]), .IN2(n5977), .Q(n47) );
  AND2X4 U232 ( .IN1(dataIn[1]), .IN2(n5978), .Q(n48) );
  AND2X4 U233 ( .IN1(dataIn[0]), .IN2(n5977), .Q(n49) );
  AND2X4 U234 ( .IN1(dataIn[8]), .IN2(n5977), .Q(n50) );
  AND2X4 U235 ( .IN1(dataIn[20]), .IN2(n5977), .Q(n51) );
  OR2X4 U236 ( .IN1(wren), .IN2(n5973), .Q(n52) );
  NBUFFX2 U237 ( .INP(n339), .Z(n6263) );
  NBUFFX2 U238 ( .INP(n339), .Z(n6262) );
  NBUFFX2 U239 ( .INP(n339), .Z(n6261) );
  NBUFFX2 U240 ( .INP(n341), .Z(n6257) );
  NBUFFX2 U241 ( .INP(n341), .Z(n6256) );
  NBUFFX2 U242 ( .INP(n341), .Z(n6255) );
  NBUFFX2 U243 ( .INP(n344), .Z(n6239) );
  NBUFFX2 U244 ( .INP(n344), .Z(n6238) );
  NBUFFX2 U245 ( .INP(n345), .Z(n6233) );
  NBUFFX2 U246 ( .INP(n345), .Z(n6232) );
  NBUFFX2 U247 ( .INP(n345), .Z(n6231) );
  NBUFFX2 U248 ( .INP(n348), .Z(n6215) );
  NBUFFX2 U249 ( .INP(n348), .Z(n6214) );
  NBUFFX2 U250 ( .INP(n349), .Z(n6209) );
  NBUFFX2 U251 ( .INP(n349), .Z(n6208) );
  NBUFFX2 U252 ( .INP(n352), .Z(n6191) );
  NBUFFX2 U253 ( .INP(n352), .Z(n6190) );
  NBUFFX2 U254 ( .INP(n352), .Z(n6189) );
  NBUFFX2 U255 ( .INP(n353), .Z(n6185) );
  NBUFFX2 U256 ( .INP(n353), .Z(n6184) );
  NBUFFX2 U257 ( .INP(n271), .Z(n6647) );
  NBUFFX2 U258 ( .INP(n271), .Z(n6646) );
  NBUFFX2 U259 ( .INP(n271), .Z(n6645) );
  NBUFFX2 U260 ( .INP(n273), .Z(n6641) );
  NBUFFX2 U261 ( .INP(n273), .Z(n6640) );
  NBUFFX2 U262 ( .INP(n273), .Z(n6639) );
  NBUFFX2 U263 ( .INP(n276), .Z(n6623) );
  NBUFFX2 U264 ( .INP(n276), .Z(n6622) );
  NBUFFX2 U265 ( .INP(n277), .Z(n6617) );
  NBUFFX2 U266 ( .INP(n277), .Z(n6616) );
  NBUFFX2 U267 ( .INP(n277), .Z(n6615) );
  NBUFFX2 U268 ( .INP(n280), .Z(n6599) );
  NBUFFX2 U269 ( .INP(n280), .Z(n6598) );
  NBUFFX2 U270 ( .INP(n281), .Z(n6593) );
  NBUFFX2 U271 ( .INP(n281), .Z(n6592) );
  NBUFFX2 U272 ( .INP(n284), .Z(n6575) );
  NBUFFX2 U273 ( .INP(n284), .Z(n6574) );
  NBUFFX2 U274 ( .INP(n284), .Z(n6573) );
  NBUFFX2 U275 ( .INP(n285), .Z(n6569) );
  NBUFFX2 U276 ( .INP(n285), .Z(n6568) );
  NBUFFX2 U277 ( .INP(n288), .Z(n6551) );
  NBUFFX2 U278 ( .INP(n288), .Z(n6550) );
  NBUFFX2 U279 ( .INP(n288), .Z(n6549) );
  NBUFFX2 U280 ( .INP(n290), .Z(n6545) );
  NBUFFX2 U281 ( .INP(n290), .Z(n6544) );
  NBUFFX2 U282 ( .INP(n293), .Z(n6527) );
  NBUFFX2 U283 ( .INP(n293), .Z(n6526) );
  NBUFFX2 U284 ( .INP(n293), .Z(n6525) );
  NBUFFX2 U285 ( .INP(n294), .Z(n6521) );
  NBUFFX2 U286 ( .INP(n294), .Z(n6520) );
  NBUFFX2 U287 ( .INP(n294), .Z(n6519) );
  NBUFFX2 U288 ( .INP(n297), .Z(n6503) );
  NBUFFX2 U289 ( .INP(n297), .Z(n6502) );
  NBUFFX2 U290 ( .INP(n297), .Z(n6501) );
  NBUFFX2 U291 ( .INP(n298), .Z(n6497) );
  NBUFFX2 U292 ( .INP(n298), .Z(n6496) );
  NBUFFX2 U293 ( .INP(n298), .Z(n6495) );
  NBUFFX2 U294 ( .INP(n301), .Z(n6479) );
  NBUFFX2 U295 ( .INP(n301), .Z(n6478) );
  NBUFFX2 U296 ( .INP(n302), .Z(n6473) );
  NBUFFX2 U297 ( .INP(n302), .Z(n6472) );
  NBUFFX2 U298 ( .INP(n302), .Z(n6471) );
  NBUFFX2 U299 ( .INP(n305), .Z(n6455) );
  NBUFFX2 U300 ( .INP(n305), .Z(n6454) );
  NBUFFX2 U301 ( .INP(n305), .Z(n6453) );
  NBUFFX2 U302 ( .INP(n307), .Z(n6449) );
  NBUFFX2 U303 ( .INP(n307), .Z(n6448) );
  NBUFFX2 U304 ( .INP(n307), .Z(n6447) );
  NBUFFX2 U305 ( .INP(n310), .Z(n6431) );
  NBUFFX2 U315 ( .INP(n310), .Z(n6430) );
  NBUFFX2 U316 ( .INP(n310), .Z(n6429) );
  NBUFFX2 U317 ( .INP(n311), .Z(n6425) );
  NBUFFX2 U318 ( .INP(n311), .Z(n6424) );
  NBUFFX2 U319 ( .INP(n311), .Z(n6423) );
  NBUFFX2 U320 ( .INP(n314), .Z(n6407) );
  NBUFFX2 U321 ( .INP(n314), .Z(n6406) );
  NBUFFX2 U322 ( .INP(n315), .Z(n6401) );
  NBUFFX2 U323 ( .INP(n315), .Z(n6400) );
  NBUFFX2 U324 ( .INP(n315), .Z(n6399) );
  NBUFFX2 U325 ( .INP(n318), .Z(n6383) );
  NBUFFX2 U326 ( .INP(n318), .Z(n6382) );
  NBUFFX2 U327 ( .INP(n319), .Z(n6377) );
  NBUFFX2 U328 ( .INP(n319), .Z(n6376) );
  NBUFFX2 U329 ( .INP(n322), .Z(n6359) );
  NBUFFX2 U330 ( .INP(n322), .Z(n6358) );
  NBUFFX2 U331 ( .INP(n324), .Z(n6353) );
  NBUFFX2 U332 ( .INP(n324), .Z(n6352) );
  NBUFFX2 U333 ( .INP(n327), .Z(n6335) );
  NBUFFX2 U334 ( .INP(n327), .Z(n6334) );
  NBUFFX2 U335 ( .INP(n327), .Z(n6333) );
  NBUFFX2 U336 ( .INP(n328), .Z(n6329) );
  NBUFFX2 U337 ( .INP(n328), .Z(n6328) );
  NBUFFX2 U338 ( .INP(n331), .Z(n6311) );
  NBUFFX2 U348 ( .INP(n331), .Z(n6310) );
  NBUFFX2 U349 ( .INP(n331), .Z(n6309) );
  NBUFFX2 U350 ( .INP(n332), .Z(n6305) );
  NBUFFX2 U351 ( .INP(n332), .Z(n6304) );
  NBUFFX2 U352 ( .INP(n332), .Z(n6303) );
  NBUFFX2 U353 ( .INP(n335), .Z(n6287) );
  NBUFFX2 U354 ( .INP(n335), .Z(n6286) );
  NBUFFX2 U355 ( .INP(n335), .Z(n6285) );
  NBUFFX2 U356 ( .INP(n336), .Z(n6281) );
  NBUFFX2 U357 ( .INP(n336), .Z(n6280) );
  NBUFFX2 U358 ( .INP(n336), .Z(n6279) );
  NBUFFX2 U359 ( .INP(n356), .Z(n6167) );
  NBUFFX2 U360 ( .INP(n356), .Z(n6166) );
  NBUFFX2 U361 ( .INP(n358), .Z(n6161) );
  NBUFFX2 U362 ( .INP(n358), .Z(n6160) );
  NBUFFX2 U363 ( .INP(n358), .Z(n6159) );
  NBUFFX2 U364 ( .INP(n361), .Z(n6143) );
  NBUFFX2 U365 ( .INP(n361), .Z(n6142) );
  NBUFFX2 U366 ( .INP(n362), .Z(n6137) );
  NBUFFX2 U367 ( .INP(n362), .Z(n6136) );
  NBUFFX2 U368 ( .INP(n365), .Z(n6119) );
  NBUFFX2 U369 ( .INP(n365), .Z(n6118) );
  NBUFFX2 U370 ( .INP(n365), .Z(n6117) );
  NBUFFX2 U371 ( .INP(n366), .Z(n6113) );
  NBUFFX2 U381 ( .INP(n366), .Z(n6112) );
  NBUFFX2 U382 ( .INP(n369), .Z(n6095) );
  NBUFFX2 U383 ( .INP(n369), .Z(n6094) );
  NBUFFX2 U384 ( .INP(n369), .Z(n6093) );
  NBUFFX2 U385 ( .INP(n370), .Z(n6089) );
  NBUFFX2 U386 ( .INP(n370), .Z(n6088) );
  NBUFFX2 U387 ( .INP(n370), .Z(n6087) );
  NBUFFX2 U388 ( .INP(n388), .Z(n6023) );
  NBUFFX2 U389 ( .INP(n388), .Z(n6022) );
  NBUFFX2 U390 ( .INP(n393), .Z(n5999) );
  NBUFFX2 U391 ( .INP(n393), .Z(n5998) );
  NBUFFX2 U392 ( .INP(n395), .Z(n5993) );
  NBUFFX2 U399 ( .INP(n395), .Z(n5992) );
  NBUFFX2 U400 ( .INP(n206), .Z(n7084) );
  NBUFFX2 U401 ( .INP(n206), .Z(n7083) );
  NBUFFX2 U402 ( .INP(n206), .Z(n7082) );
  NBUFFX2 U403 ( .INP(n240), .Z(n6737) );
  NBUFFX2 U404 ( .INP(n240), .Z(n6736) );
  NBUFFX2 U414 ( .INP(n240), .Z(n6735) );
  NBUFFX2 U415 ( .INP(n242), .Z(n6731) );
  NBUFFX2 U416 ( .INP(n242), .Z(n6730) );
  NBUFFX2 U417 ( .INP(n244), .Z(n6725) );
  NBUFFX2 U418 ( .INP(n246), .Z(n6719) );
  NBUFFX2 U419 ( .INP(n246), .Z(n6718) );
  NBUFFX2 U420 ( .INP(n246), .Z(n6717) );
  NBUFFX2 U421 ( .INP(n248), .Z(n6713) );
  NBUFFX2 U422 ( .INP(n248), .Z(n6712) );
  NBUFFX2 U423 ( .INP(n248), .Z(n6711) );
  NBUFFX2 U424 ( .INP(n254), .Z(n6695) );
  NBUFFX2 U425 ( .INP(n254), .Z(n6694) );
  NBUFFX2 U426 ( .INP(n256), .Z(n6689) );
  NBUFFX2 U427 ( .INP(n256), .Z(n6688) );
  NBUFFX2 U428 ( .INP(n256), .Z(n6687) );
  NBUFFX2 U429 ( .INP(n262), .Z(n6671) );
  NBUFFX2 U430 ( .INP(n262), .Z(n6670) );
  NBUFFX2 U431 ( .INP(n264), .Z(n6665) );
  NBUFFX2 U432 ( .INP(n264), .Z(n6664) );
  NBUFFX2 U433 ( .INP(n244), .Z(n6724) );
  NBUFFX2 U434 ( .INP(n344), .Z(n6237) );
  NBUFFX2 U435 ( .INP(n348), .Z(n6213) );
  NBUFFX2 U436 ( .INP(n349), .Z(n6207) );
  NBUFFX2 U437 ( .INP(n353), .Z(n6183) );
  NBUFFX2 U447 ( .INP(n276), .Z(n6621) );
  NBUFFX2 U448 ( .INP(n280), .Z(n6597) );
  NBUFFX2 U449 ( .INP(n281), .Z(n6591) );
  NBUFFX2 U450 ( .INP(n285), .Z(n6567) );
  NBUFFX2 U451 ( .INP(n290), .Z(n6543) );
  NBUFFX2 U452 ( .INP(n301), .Z(n6477) );
  NBUFFX2 U453 ( .INP(n314), .Z(n6405) );
  NBUFFX2 U454 ( .INP(n318), .Z(n6381) );
  NBUFFX2 U455 ( .INP(n319), .Z(n6375) );
  NBUFFX2 U456 ( .INP(n322), .Z(n6357) );
  NBUFFX2 U457 ( .INP(n324), .Z(n6351) );
  NBUFFX2 U458 ( .INP(n328), .Z(n6327) );
  NBUFFX2 U459 ( .INP(n356), .Z(n6165) );
  NBUFFX2 U460 ( .INP(n361), .Z(n6141) );
  NBUFFX2 U461 ( .INP(n362), .Z(n6135) );
  NBUFFX2 U462 ( .INP(n366), .Z(n6111) );
  NBUFFX2 U463 ( .INP(n388), .Z(n6021) );
  NBUFFX2 U464 ( .INP(n393), .Z(n5997) );
  NBUFFX2 U465 ( .INP(n395), .Z(n5991) );
  NBUFFX2 U466 ( .INP(n242), .Z(n6729) );
  NBUFFX2 U467 ( .INP(n244), .Z(n6723) );
  NBUFFX2 U468 ( .INP(n254), .Z(n6693) );
  NBUFFX2 U469 ( .INP(n262), .Z(n6669) );
  NBUFFX2 U470 ( .INP(n264), .Z(n6663) );
  NBUFFX2 U546 ( .INP(n342), .Z(n6251) );
  NBUFFX2 U547 ( .INP(n342), .Z(n6250) );
  NBUFFX2 U548 ( .INP(n342), .Z(n6249) );
  NBUFFX2 U549 ( .INP(n343), .Z(n6245) );
  NBUFFX2 U550 ( .INP(n343), .Z(n6244) );
  NBUFFX2 U551 ( .INP(n343), .Z(n6243) );
  NBUFFX2 U552 ( .INP(n346), .Z(n6227) );
  NBUFFX2 U553 ( .INP(n346), .Z(n6226) );
  NBUFFX2 U554 ( .INP(n346), .Z(n6225) );
  NBUFFX2 U555 ( .INP(n347), .Z(n6221) );
  NBUFFX2 U556 ( .INP(n347), .Z(n6220) );
  NBUFFX2 U557 ( .INP(n347), .Z(n6219) );
  NBUFFX2 U558 ( .INP(n350), .Z(n6203) );
  NBUFFX2 U559 ( .INP(n350), .Z(n6202) );
  NBUFFX2 U560 ( .INP(n350), .Z(n6201) );
  NBUFFX2 U561 ( .INP(n351), .Z(n6197) );
  NBUFFX2 U562 ( .INP(n351), .Z(n6196) );
  NBUFFX2 U563 ( .INP(n351), .Z(n6195) );
  NBUFFX2 U564 ( .INP(n354), .Z(n6179) );
  NBUFFX2 U565 ( .INP(n354), .Z(n6178) );
  NBUFFX2 U566 ( .INP(n354), .Z(n6177) );
  NBUFFX2 U567 ( .INP(n355), .Z(n6173) );
  NBUFFX2 U568 ( .INP(n355), .Z(n6172) );
  NBUFFX2 U569 ( .INP(n355), .Z(n6171) );
  NBUFFX2 U579 ( .INP(n250), .Z(n6707) );
  NBUFFX2 U580 ( .INP(n250), .Z(n6706) );
  NBUFFX2 U581 ( .INP(n250), .Z(n6705) );
  NBUFFX2 U582 ( .INP(n252), .Z(n6701) );
  NBUFFX2 U583 ( .INP(n252), .Z(n6700) );
  NBUFFX2 U584 ( .INP(n252), .Z(n6699) );
  NBUFFX2 U585 ( .INP(n258), .Z(n6683) );
  NBUFFX2 U586 ( .INP(n258), .Z(n6682) );
  NBUFFX2 U587 ( .INP(n258), .Z(n6681) );
  NBUFFX2 U588 ( .INP(n260), .Z(n6677) );
  NBUFFX2 U589 ( .INP(n260), .Z(n6676) );
  NBUFFX2 U590 ( .INP(n260), .Z(n6675) );
  NBUFFX2 U591 ( .INP(n266), .Z(n6659) );
  NBUFFX2 U592 ( .INP(n266), .Z(n6658) );
  NBUFFX2 U593 ( .INP(n266), .Z(n6657) );
  NBUFFX2 U594 ( .INP(n268), .Z(n6653) );
  NBUFFX2 U595 ( .INP(n268), .Z(n6652) );
  NBUFFX2 U596 ( .INP(n268), .Z(n6651) );
  NBUFFX2 U597 ( .INP(n274), .Z(n6635) );
  NBUFFX2 U598 ( .INP(n274), .Z(n6634) );
  NBUFFX2 U599 ( .INP(n274), .Z(n6633) );
  NBUFFX2 U600 ( .INP(n275), .Z(n6629) );
  NBUFFX2 U601 ( .INP(n275), .Z(n6628) );
  NBUFFX2 U602 ( .INP(n275), .Z(n6627) );
  NBUFFX2 U678 ( .INP(n278), .Z(n6611) );
  NBUFFX2 U679 ( .INP(n278), .Z(n6610) );
  NBUFFX2 U680 ( .INP(n278), .Z(n6609) );
  NBUFFX2 U681 ( .INP(n279), .Z(n6605) );
  NBUFFX2 U682 ( .INP(n279), .Z(n6604) );
  NBUFFX2 U683 ( .INP(n279), .Z(n6603) );
  NBUFFX2 U684 ( .INP(n282), .Z(n6587) );
  NBUFFX2 U685 ( .INP(n282), .Z(n6586) );
  NBUFFX2 U686 ( .INP(n282), .Z(n6585) );
  NBUFFX2 U687 ( .INP(n283), .Z(n6581) );
  NBUFFX2 U688 ( .INP(n283), .Z(n6580) );
  NBUFFX2 U689 ( .INP(n283), .Z(n6579) );
  NBUFFX2 U690 ( .INP(n286), .Z(n6563) );
  NBUFFX2 U691 ( .INP(n286), .Z(n6562) );
  NBUFFX2 U692 ( .INP(n286), .Z(n6561) );
  NBUFFX2 U693 ( .INP(n287), .Z(n6557) );
  NBUFFX2 U694 ( .INP(n287), .Z(n6556) );
  NBUFFX2 U695 ( .INP(n287), .Z(n6555) );
  NBUFFX2 U696 ( .INP(n291), .Z(n6539) );
  NBUFFX2 U697 ( .INP(n291), .Z(n6538) );
  NBUFFX2 U698 ( .INP(n291), .Z(n6537) );
  NBUFFX2 U699 ( .INP(n292), .Z(n6533) );
  NBUFFX2 U700 ( .INP(n292), .Z(n6532) );
  NBUFFX2 U701 ( .INP(n292), .Z(n6531) );
  NBUFFX2 U711 ( .INP(n295), .Z(n6515) );
  NBUFFX2 U712 ( .INP(n295), .Z(n6514) );
  NBUFFX2 U713 ( .INP(n295), .Z(n6513) );
  NBUFFX2 U714 ( .INP(n296), .Z(n6509) );
  NBUFFX2 U715 ( .INP(n296), .Z(n6508) );
  NBUFFX2 U716 ( .INP(n296), .Z(n6507) );
  NBUFFX2 U717 ( .INP(n299), .Z(n6491) );
  NBUFFX2 U718 ( .INP(n299), .Z(n6490) );
  NBUFFX2 U719 ( .INP(n299), .Z(n6489) );
  NBUFFX2 U720 ( .INP(n300), .Z(n6485) );
  NBUFFX2 U721 ( .INP(n300), .Z(n6484) );
  NBUFFX2 U722 ( .INP(n300), .Z(n6483) );
  NBUFFX2 U723 ( .INP(n303), .Z(n6467) );
  NBUFFX2 U724 ( .INP(n303), .Z(n6466) );
  NBUFFX2 U725 ( .INP(n303), .Z(n6465) );
  NBUFFX2 U726 ( .INP(n304), .Z(n6461) );
  NBUFFX2 U727 ( .INP(n304), .Z(n6460) );
  NBUFFX2 U728 ( .INP(n304), .Z(n6459) );
  NBUFFX2 U729 ( .INP(n308), .Z(n6443) );
  NBUFFX2 U730 ( .INP(n308), .Z(n6442) );
  NBUFFX2 U731 ( .INP(n308), .Z(n6441) );
  NBUFFX2 U732 ( .INP(n309), .Z(n6437) );
  NBUFFX2 U733 ( .INP(n309), .Z(n6436) );
  NBUFFX2 U734 ( .INP(n309), .Z(n6435) );
  NBUFFX2 U751 ( .INP(n312), .Z(n6419) );
  NBUFFX2 U810 ( .INP(n312), .Z(n6418) );
  NBUFFX2 U811 ( .INP(n312), .Z(n6417) );
  NBUFFX2 U812 ( .INP(n313), .Z(n6413) );
  NBUFFX2 U813 ( .INP(n313), .Z(n6412) );
  NBUFFX2 U814 ( .INP(n313), .Z(n6411) );
  NBUFFX2 U815 ( .INP(n316), .Z(n6395) );
  NBUFFX2 U816 ( .INP(n316), .Z(n6394) );
  NBUFFX2 U817 ( .INP(n316), .Z(n6393) );
  NBUFFX2 U818 ( .INP(n317), .Z(n6389) );
  NBUFFX2 U819 ( .INP(n317), .Z(n6388) );
  NBUFFX2 U820 ( .INP(n317), .Z(n6387) );
  NBUFFX2 U821 ( .INP(n320), .Z(n6371) );
  NBUFFX2 U822 ( .INP(n320), .Z(n6370) );
  NBUFFX2 U823 ( .INP(n320), .Z(n6369) );
  NBUFFX2 U824 ( .INP(n321), .Z(n6365) );
  NBUFFX2 U825 ( .INP(n321), .Z(n6364) );
  NBUFFX2 U826 ( .INP(n321), .Z(n6363) );
  NBUFFX2 U827 ( .INP(n325), .Z(n6347) );
  NBUFFX2 U828 ( .INP(n325), .Z(n6346) );
  NBUFFX2 U829 ( .INP(n325), .Z(n6345) );
  NBUFFX2 U830 ( .INP(n326), .Z(n6341) );
  NBUFFX2 U831 ( .INP(n326), .Z(n6340) );
  NBUFFX2 U832 ( .INP(n326), .Z(n6339) );
  NBUFFX2 U833 ( .INP(n329), .Z(n6323) );
  NBUFFX2 U834 ( .INP(n329), .Z(n6322) );
  NBUFFX2 U844 ( .INP(n329), .Z(n6321) );
  NBUFFX2 U845 ( .INP(n330), .Z(n6317) );
  NBUFFX2 U846 ( .INP(n330), .Z(n6316) );
  NBUFFX2 U847 ( .INP(n330), .Z(n6315) );
  NBUFFX2 U848 ( .INP(n333), .Z(n6299) );
  NBUFFX2 U849 ( .INP(n333), .Z(n6298) );
  NBUFFX2 U850 ( .INP(n333), .Z(n6297) );
  NBUFFX2 U851 ( .INP(n334), .Z(n6293) );
  NBUFFX2 U852 ( .INP(n334), .Z(n6292) );
  NBUFFX2 U853 ( .INP(n334), .Z(n6291) );
  NBUFFX2 U854 ( .INP(n337), .Z(n6275) );
  NBUFFX2 U855 ( .INP(n337), .Z(n6274) );
  NBUFFX2 U856 ( .INP(n337), .Z(n6273) );
  NBUFFX2 U857 ( .INP(n338), .Z(n6269) );
  NBUFFX2 U858 ( .INP(n338), .Z(n6268) );
  NBUFFX2 U859 ( .INP(n338), .Z(n6267) );
  NBUFFX2 U860 ( .INP(n359), .Z(n6155) );
  NBUFFX2 U861 ( .INP(n359), .Z(n6154) );
  NBUFFX2 U862 ( .INP(n359), .Z(n6153) );
  NBUFFX2 U863 ( .INP(n360), .Z(n6149) );
  NBUFFX2 U864 ( .INP(n360), .Z(n6148) );
  NBUFFX2 U865 ( .INP(n360), .Z(n6147) );
  NBUFFX2 U866 ( .INP(n363), .Z(n6131) );
  NBUFFX2 U867 ( .INP(n363), .Z(n6130) );
  NBUFFX2 U918 ( .INP(n363), .Z(n6129) );
  NBUFFX2 U943 ( .INP(n364), .Z(n6125) );
  NBUFFX2 U944 ( .INP(n364), .Z(n6124) );
  NBUFFX2 U945 ( .INP(n364), .Z(n6123) );
  NBUFFX2 U946 ( .INP(n367), .Z(n6107) );
  NBUFFX2 U947 ( .INP(n367), .Z(n6106) );
  NBUFFX2 U948 ( .INP(n367), .Z(n6105) );
  NBUFFX2 U949 ( .INP(n368), .Z(n6101) );
  NBUFFX2 U950 ( .INP(n368), .Z(n6100) );
  NBUFFX2 U951 ( .INP(n368), .Z(n6099) );
  NBUFFX2 U952 ( .INP(n371), .Z(n6083) );
  NBUFFX2 U953 ( .INP(n371), .Z(n6082) );
  NBUFFX2 U954 ( .INP(n371), .Z(n6081) );
  NBUFFX2 U955 ( .INP(n372), .Z(n6077) );
  NBUFFX2 U956 ( .INP(n372), .Z(n6076) );
  NBUFFX2 U957 ( .INP(n372), .Z(n6075) );
  NBUFFX2 U958 ( .INP(n379), .Z(n6059) );
  NBUFFX2 U959 ( .INP(n379), .Z(n6058) );
  NBUFFX2 U960 ( .INP(n379), .Z(n6057) );
  NBUFFX2 U961 ( .INP(n381), .Z(n6053) );
  NBUFFX2 U962 ( .INP(n381), .Z(n6052) );
  NBUFFX2 U963 ( .INP(n381), .Z(n6051) );
  NBUFFX2 U964 ( .INP(n387), .Z(n6029) );
  NBUFFX2 U965 ( .INP(n387), .Z(n6028) );
  NBUFFX2 U966 ( .INP(n387), .Z(n6027) );
  NBUFFX2 U976 ( .INP(n392), .Z(n6005) );
  NBUFFX2 U977 ( .INP(n392), .Z(n6004) );
  NBUFFX2 U978 ( .INP(n392), .Z(n6003) );
  NBUFFX2 U979 ( .INP(n396), .Z(n5987) );
  NBUFFX2 U980 ( .INP(n396), .Z(n5986) );
  NBUFFX2 U981 ( .INP(n396), .Z(n5985) );
  NBUFFX2 U982 ( .INP(n397), .Z(n5981) );
  NBUFFX2 U983 ( .INP(n397), .Z(n5980) );
  NBUFFX2 U984 ( .INP(n397), .Z(n5979) );
  NBUFFX2 U985 ( .INP(n7357), .Z(n7334) );
  NBUFFX2 U986 ( .INP(n7357), .Z(n7335) );
  NBUFFX2 U987 ( .INP(n7357), .Z(n7336) );
  NBUFFX2 U988 ( .INP(n7356), .Z(n7337) );
  NBUFFX2 U989 ( .INP(n7356), .Z(n7338) );
  NBUFFX2 U990 ( .INP(n7356), .Z(n7339) );
  NBUFFX2 U991 ( .INP(n7344), .Z(n7340) );
  NBUFFX2 U992 ( .INP(n7355), .Z(n7341) );
  NBUFFX2 U993 ( .INP(n7355), .Z(n7342) );
  NBUFFX2 U994 ( .INP(n7355), .Z(n7343) );
  NBUFFX2 U995 ( .INP(n7351), .Z(n7344) );
  NBUFFX2 U996 ( .INP(n7352), .Z(n7345) );
  NBUFFX2 U997 ( .INP(n7347), .Z(n7346) );
  NBUFFX2 U998 ( .INP(n7354), .Z(n7347) );
  NBUFFX2 U999 ( .INP(n7354), .Z(n7348) );
  NBUFFX2 U1075 ( .INP(n7354), .Z(n7349) );
  NBUFFX2 U1076 ( .INP(n7353), .Z(n7350) );
  NBUFFX2 U1077 ( .INP(n7353), .Z(n7351) );
  NBUFFX2 U1078 ( .INP(n7353), .Z(n7352) );
  NOR2X0 U1079 ( .IN1(n7363), .IN2(n7362), .QN(n376) );
  NOR2X0 U1080 ( .IN1(n7365), .IN2(n7364), .QN(n375) );
  NBUFFX2 U1081 ( .INP(n49), .Z(n7097) );
  NBUFFX2 U1082 ( .INP(n48), .Z(n7080) );
  NBUFFX2 U1083 ( .INP(n47), .Z(n7069) );
  NBUFFX2 U1084 ( .INP(n46), .Z(n7058) );
  NBUFFX2 U1085 ( .INP(n45), .Z(n7047) );
  NBUFFX2 U1086 ( .INP(n44), .Z(n7036) );
  NBUFFX2 U1087 ( .INP(n43), .Z(n7025) );
  NBUFFX2 U1088 ( .INP(n42), .Z(n7014) );
  NBUFFX2 U1089 ( .INP(n50), .Z(n7003) );
  NBUFFX2 U1090 ( .INP(n27), .Z(n6992) );
  NBUFFX2 U1091 ( .INP(n26), .Z(n6981) );
  NBUFFX2 U1092 ( .INP(n25), .Z(n6970) );
  NBUFFX2 U1093 ( .INP(n33), .Z(n6959) );
  NBUFFX2 U1094 ( .INP(n32), .Z(n6948) );
  NBUFFX2 U1095 ( .INP(n31), .Z(n6937) );
  NBUFFX2 U1096 ( .INP(n30), .Z(n6926) );
  NBUFFX2 U1097 ( .INP(n29), .Z(n6915) );
  NBUFFX2 U1098 ( .INP(n28), .Z(n6904) );
  NBUFFX2 U1108 ( .INP(n24), .Z(n6893) );
  NBUFFX2 U1109 ( .INP(n23), .Z(n6882) );
  NBUFFX2 U1110 ( .INP(n51), .Z(n6871) );
  NBUFFX2 U1111 ( .INP(n22), .Z(n6860) );
  NBUFFX2 U1112 ( .INP(n21), .Z(n6849) );
  NBUFFX2 U1113 ( .INP(n20), .Z(n6838) );
  NBUFFX2 U1114 ( .INP(n49), .Z(n7096) );
  NBUFFX2 U1115 ( .INP(n48), .Z(n7079) );
  NBUFFX2 U1116 ( .INP(n47), .Z(n7068) );
  NBUFFX2 U1117 ( .INP(n46), .Z(n7057) );
  NBUFFX2 U1118 ( .INP(n45), .Z(n7046) );
  NBUFFX2 U1119 ( .INP(n44), .Z(n7035) );
  NBUFFX2 U1120 ( .INP(n43), .Z(n7024) );
  NBUFFX2 U1121 ( .INP(n42), .Z(n7013) );
  NBUFFX2 U1122 ( .INP(n50), .Z(n7002) );
  NBUFFX2 U1123 ( .INP(n27), .Z(n6991) );
  NBUFFX2 U1124 ( .INP(n26), .Z(n6980) );
  NBUFFX2 U1125 ( .INP(n25), .Z(n6969) );
  NBUFFX2 U1126 ( .INP(n33), .Z(n6958) );
  NBUFFX2 U1127 ( .INP(n32), .Z(n6947) );
  NBUFFX2 U1128 ( .INP(n31), .Z(n6936) );
  NBUFFX2 U1129 ( .INP(n30), .Z(n6925) );
  NBUFFX2 U1130 ( .INP(n29), .Z(n6914) );
  NBUFFX2 U1131 ( .INP(n28), .Z(n6903) );
  NBUFFX2 U1207 ( .INP(n24), .Z(n6892) );
  NBUFFX2 U1208 ( .INP(n23), .Z(n6881) );
  NBUFFX2 U1209 ( .INP(n51), .Z(n6870) );
  NBUFFX2 U1210 ( .INP(n22), .Z(n6859) );
  NBUFFX2 U1211 ( .INP(n21), .Z(n6848) );
  NBUFFX2 U1212 ( .INP(n20), .Z(n6837) );
  NBUFFX2 U1213 ( .INP(n49), .Z(n7095) );
  NBUFFX2 U1214 ( .INP(n48), .Z(n7078) );
  NBUFFX2 U1215 ( .INP(n47), .Z(n7067) );
  NBUFFX2 U1216 ( .INP(n46), .Z(n7056) );
  NBUFFX2 U1217 ( .INP(n45), .Z(n7045) );
  NBUFFX2 U1218 ( .INP(n44), .Z(n7034) );
  NBUFFX2 U1219 ( .INP(n43), .Z(n7023) );
  NBUFFX2 U1220 ( .INP(n42), .Z(n7012) );
  NBUFFX2 U1221 ( .INP(n50), .Z(n7001) );
  NBUFFX2 U1222 ( .INP(n27), .Z(n6990) );
  NBUFFX2 U1223 ( .INP(n26), .Z(n6979) );
  NBUFFX2 U1224 ( .INP(n25), .Z(n6968) );
  NBUFFX2 U1225 ( .INP(n33), .Z(n6957) );
  NBUFFX2 U1226 ( .INP(n32), .Z(n6946) );
  NBUFFX2 U1227 ( .INP(n31), .Z(n6935) );
  NBUFFX2 U1228 ( .INP(n30), .Z(n6924) );
  NBUFFX2 U1229 ( .INP(n29), .Z(n6913) );
  NBUFFX2 U1230 ( .INP(n28), .Z(n6902) );
  NBUFFX2 U1240 ( .INP(n24), .Z(n6891) );
  NBUFFX2 U1241 ( .INP(n23), .Z(n6880) );
  NBUFFX2 U1242 ( .INP(n51), .Z(n6869) );
  NBUFFX2 U1243 ( .INP(n22), .Z(n6858) );
  NBUFFX2 U1244 ( .INP(n21), .Z(n6847) );
  NBUFFX2 U1245 ( .INP(n20), .Z(n6836) );
  NBUFFX2 U1246 ( .INP(n49), .Z(n7094) );
  NBUFFX2 U1247 ( .INP(n48), .Z(n7077) );
  NBUFFX2 U1248 ( .INP(n47), .Z(n7066) );
  NBUFFX2 U1249 ( .INP(n46), .Z(n7055) );
  NBUFFX2 U1250 ( .INP(n45), .Z(n7044) );
  NBUFFX2 U1251 ( .INP(n44), .Z(n7033) );
  NBUFFX2 U1252 ( .INP(n43), .Z(n7022) );
  NBUFFX2 U1253 ( .INP(n42), .Z(n7011) );
  NBUFFX2 U1254 ( .INP(n50), .Z(n7000) );
  NBUFFX2 U1255 ( .INP(n27), .Z(n6989) );
  NBUFFX2 U1256 ( .INP(n26), .Z(n6978) );
  NBUFFX2 U1257 ( .INP(n25), .Z(n6967) );
  NBUFFX2 U1258 ( .INP(n33), .Z(n6956) );
  NBUFFX2 U1259 ( .INP(n32), .Z(n6945) );
  NBUFFX2 U1260 ( .INP(n31), .Z(n6934) );
  NBUFFX2 U1261 ( .INP(n30), .Z(n6923) );
  NBUFFX2 U1262 ( .INP(n29), .Z(n6912) );
  NBUFFX2 U1263 ( .INP(n28), .Z(n6901) );
  NBUFFX2 U1273 ( .INP(n24), .Z(n6890) );
  NBUFFX2 U1287 ( .INP(n23), .Z(n6879) );
  NBUFFX2 U1339 ( .INP(n51), .Z(n6868) );
  NBUFFX2 U1340 ( .INP(n22), .Z(n6857) );
  NBUFFX2 U1341 ( .INP(n21), .Z(n6846) );
  NBUFFX2 U1342 ( .INP(n20), .Z(n6835) );
  NBUFFX2 U1343 ( .INP(n49), .Z(n7093) );
  NBUFFX2 U1344 ( .INP(n48), .Z(n7076) );
  NBUFFX2 U1345 ( .INP(n47), .Z(n7065) );
  NBUFFX2 U1346 ( .INP(n46), .Z(n7054) );
  NBUFFX2 U1347 ( .INP(n45), .Z(n7043) );
  NBUFFX2 U1348 ( .INP(n44), .Z(n7032) );
  NBUFFX2 U1349 ( .INP(n43), .Z(n7021) );
  NBUFFX2 U1350 ( .INP(n42), .Z(n7010) );
  NBUFFX2 U1351 ( .INP(n50), .Z(n6999) );
  NBUFFX2 U1352 ( .INP(n27), .Z(n6988) );
  NBUFFX2 U1353 ( .INP(n26), .Z(n6977) );
  NBUFFX2 U1354 ( .INP(n25), .Z(n6966) );
  NBUFFX2 U1355 ( .INP(n33), .Z(n6955) );
  NBUFFX2 U1356 ( .INP(n32), .Z(n6944) );
  NBUFFX2 U1357 ( .INP(n31), .Z(n6933) );
  NBUFFX2 U1358 ( .INP(n30), .Z(n6922) );
  NBUFFX2 U1359 ( .INP(n29), .Z(n6911) );
  NBUFFX2 U1360 ( .INP(n28), .Z(n6900) );
  NBUFFX2 U1361 ( .INP(n24), .Z(n6889) );
  NBUFFX2 U1362 ( .INP(n23), .Z(n6878) );
  NBUFFX2 U1363 ( .INP(n51), .Z(n6867) );
  NBUFFX2 U1373 ( .INP(n22), .Z(n6856) );
  NBUFFX2 U1374 ( .INP(n21), .Z(n6845) );
  NBUFFX2 U1375 ( .INP(n20), .Z(n6834) );
  NBUFFX2 U1376 ( .INP(n49), .Z(n7092) );
  NBUFFX2 U1377 ( .INP(n48), .Z(n7075) );
  NBUFFX2 U1378 ( .INP(n47), .Z(n7064) );
  NBUFFX2 U1379 ( .INP(n46), .Z(n7053) );
  NBUFFX2 U1380 ( .INP(n45), .Z(n7042) );
  NBUFFX2 U1381 ( .INP(n44), .Z(n7031) );
  NBUFFX2 U1382 ( .INP(n43), .Z(n7020) );
  NBUFFX2 U1383 ( .INP(n42), .Z(n7009) );
  NBUFFX2 U1384 ( .INP(n50), .Z(n6998) );
  NBUFFX2 U1385 ( .INP(n27), .Z(n6987) );
  NBUFFX2 U1386 ( .INP(n26), .Z(n6976) );
  NBUFFX2 U1387 ( .INP(n25), .Z(n6965) );
  NBUFFX2 U1388 ( .INP(n33), .Z(n6954) );
  NBUFFX2 U1389 ( .INP(n32), .Z(n6943) );
  NBUFFX2 U1390 ( .INP(n31), .Z(n6932) );
  NBUFFX2 U1391 ( .INP(n30), .Z(n6921) );
  NBUFFX2 U1392 ( .INP(n29), .Z(n6910) );
  NBUFFX2 U1393 ( .INP(n28), .Z(n6899) );
  NBUFFX2 U1394 ( .INP(n24), .Z(n6888) );
  NBUFFX2 U1395 ( .INP(n23), .Z(n6877) );
  NBUFFX2 U1396 ( .INP(n51), .Z(n6866) );
  NBUFFX2 U1408 ( .INP(n22), .Z(n6855) );
  NBUFFX2 U1423 ( .INP(n21), .Z(n6844) );
  NBUFFX2 U1472 ( .INP(n20), .Z(n6833) );
  NBUFFX2 U1473 ( .INP(n49), .Z(n7091) );
  NBUFFX2 U1474 ( .INP(n48), .Z(n7074) );
  NBUFFX2 U1475 ( .INP(n47), .Z(n7063) );
  NBUFFX2 U1476 ( .INP(n46), .Z(n7052) );
  NBUFFX2 U1477 ( .INP(n45), .Z(n7041) );
  NBUFFX2 U1478 ( .INP(n44), .Z(n7030) );
  NBUFFX2 U1479 ( .INP(n43), .Z(n7019) );
  NBUFFX2 U1480 ( .INP(n42), .Z(n7008) );
  NBUFFX2 U1481 ( .INP(n50), .Z(n6997) );
  NBUFFX2 U1482 ( .INP(n27), .Z(n6986) );
  NBUFFX2 U1483 ( .INP(n26), .Z(n6975) );
  NBUFFX2 U1484 ( .INP(n25), .Z(n6964) );
  NBUFFX2 U1485 ( .INP(n33), .Z(n6953) );
  NBUFFX2 U1486 ( .INP(n32), .Z(n6942) );
  NBUFFX2 U1487 ( .INP(n31), .Z(n6931) );
  NBUFFX2 U1488 ( .INP(n30), .Z(n6920) );
  NBUFFX2 U1489 ( .INP(n29), .Z(n6909) );
  NBUFFX2 U1490 ( .INP(n28), .Z(n6898) );
  NBUFFX2 U1491 ( .INP(n24), .Z(n6887) );
  NBUFFX2 U1492 ( .INP(n23), .Z(n6876) );
  NBUFFX2 U1493 ( .INP(n51), .Z(n6865) );
  NBUFFX2 U1494 ( .INP(n22), .Z(n6854) );
  NBUFFX2 U1495 ( .INP(n21), .Z(n6843) );
  NBUFFX2 U1505 ( .INP(n20), .Z(n6832) );
  NBUFFX2 U1506 ( .INP(n49), .Z(n7090) );
  NBUFFX2 U1507 ( .INP(n48), .Z(n7073) );
  NBUFFX2 U1508 ( .INP(n47), .Z(n7062) );
  NBUFFX2 U1509 ( .INP(n46), .Z(n7051) );
  NBUFFX2 U1510 ( .INP(n45), .Z(n7040) );
  NBUFFX2 U1511 ( .INP(n44), .Z(n7029) );
  NBUFFX2 U1512 ( .INP(n43), .Z(n7018) );
  NBUFFX2 U1513 ( .INP(n42), .Z(n7007) );
  NBUFFX2 U1514 ( .INP(n50), .Z(n6996) );
  NBUFFX2 U1515 ( .INP(n27), .Z(n6985) );
  NBUFFX2 U1516 ( .INP(n26), .Z(n6974) );
  NBUFFX2 U1517 ( .INP(n25), .Z(n6963) );
  NBUFFX2 U1518 ( .INP(n33), .Z(n6952) );
  NBUFFX2 U1519 ( .INP(n32), .Z(n6941) );
  NBUFFX2 U1520 ( .INP(n31), .Z(n6930) );
  NBUFFX2 U1521 ( .INP(n30), .Z(n6919) );
  NBUFFX2 U1522 ( .INP(n29), .Z(n6908) );
  NBUFFX2 U1523 ( .INP(n28), .Z(n6897) );
  NBUFFX2 U1524 ( .INP(n24), .Z(n6886) );
  NBUFFX2 U1525 ( .INP(n23), .Z(n6875) );
  NBUFFX2 U1526 ( .INP(n51), .Z(n6864) );
  NBUFFX2 U1527 ( .INP(n22), .Z(n6853) );
  NBUFFX2 U1528 ( .INP(n21), .Z(n6842) );
  NBUFFX2 U1541 ( .INP(n20), .Z(n6831) );
  NBUFFX2 U1554 ( .INP(n49), .Z(n7089) );
  NBUFFX2 U1575 ( .INP(n48), .Z(n7072) );
  NBUFFX2 U1604 ( .INP(n47), .Z(n7061) );
  NBUFFX2 U1605 ( .INP(n46), .Z(n7050) );
  NBUFFX2 U1606 ( .INP(n45), .Z(n7039) );
  NBUFFX2 U1607 ( .INP(n44), .Z(n7028) );
  NBUFFX2 U1608 ( .INP(n43), .Z(n7017) );
  NBUFFX2 U1609 ( .INP(n42), .Z(n7006) );
  NBUFFX2 U1610 ( .INP(n50), .Z(n6995) );
  NBUFFX2 U1611 ( .INP(n27), .Z(n6984) );
  NBUFFX2 U1612 ( .INP(n26), .Z(n6973) );
  NBUFFX2 U1613 ( .INP(n25), .Z(n6962) );
  NBUFFX2 U1614 ( .INP(n33), .Z(n6951) );
  NBUFFX2 U1615 ( .INP(n32), .Z(n6940) );
  NBUFFX2 U1616 ( .INP(n31), .Z(n6929) );
  NBUFFX2 U1617 ( .INP(n30), .Z(n6918) );
  NBUFFX2 U1618 ( .INP(n29), .Z(n6907) );
  NBUFFX2 U1619 ( .INP(n28), .Z(n6896) );
  NBUFFX2 U1620 ( .INP(n24), .Z(n6885) );
  NBUFFX2 U1621 ( .INP(n23), .Z(n6874) );
  NBUFFX2 U1622 ( .INP(n51), .Z(n6863) );
  NBUFFX2 U1623 ( .INP(n22), .Z(n6852) );
  NBUFFX2 U1624 ( .INP(n21), .Z(n6841) );
  NBUFFX2 U1625 ( .INP(n20), .Z(n6830) );
  NBUFFX2 U1626 ( .INP(n49), .Z(n7088) );
  NBUFFX2 U1627 ( .INP(n48), .Z(n7071) );
  NBUFFX2 U1637 ( .INP(n47), .Z(n7060) );
  NBUFFX2 U1638 ( .INP(n46), .Z(n7049) );
  NBUFFX2 U1639 ( .INP(n45), .Z(n7038) );
  NBUFFX2 U1640 ( .INP(n44), .Z(n7027) );
  NBUFFX2 U1641 ( .INP(n43), .Z(n7016) );
  NBUFFX2 U1642 ( .INP(n42), .Z(n7005) );
  NBUFFX2 U1643 ( .INP(n50), .Z(n6994) );
  NBUFFX2 U1644 ( .INP(n27), .Z(n6983) );
  NBUFFX2 U1645 ( .INP(n26), .Z(n6972) );
  NBUFFX2 U1646 ( .INP(n25), .Z(n6961) );
  NBUFFX2 U1647 ( .INP(n33), .Z(n6950) );
  NBUFFX2 U1648 ( .INP(n32), .Z(n6939) );
  NBUFFX2 U1649 ( .INP(n31), .Z(n6928) );
  NBUFFX2 U1650 ( .INP(n30), .Z(n6917) );
  NBUFFX2 U1651 ( .INP(n29), .Z(n6906) );
  NBUFFX2 U1652 ( .INP(n28), .Z(n6895) );
  NBUFFX2 U1653 ( .INP(n24), .Z(n6884) );
  NBUFFX2 U1654 ( .INP(n23), .Z(n6873) );
  NBUFFX2 U1655 ( .INP(n51), .Z(n6862) );
  NBUFFX2 U1656 ( .INP(n22), .Z(n6851) );
  NBUFFX2 U1657 ( .INP(n21), .Z(n6840) );
  NBUFFX2 U1658 ( .INP(n20), .Z(n6829) );
  NBUFFX2 U1659 ( .INP(n41), .Z(n6827) );
  NBUFFX2 U1660 ( .INP(n40), .Z(n6816) );
  NBUFFX2 U1708 ( .INP(n39), .Z(n6805) );
  NBUFFX2 U1721 ( .INP(n38), .Z(n6794) );
  NBUFFX2 U1736 ( .INP(n37), .Z(n6783) );
  NBUFFX2 U1737 ( .INP(n36), .Z(n6772) );
  NBUFFX2 U1738 ( .INP(n35), .Z(n6761) );
  NBUFFX2 U1739 ( .INP(n34), .Z(n6750) );
  NBUFFX2 U1740 ( .INP(n41), .Z(n6826) );
  NBUFFX2 U1741 ( .INP(n40), .Z(n6815) );
  NBUFFX2 U1742 ( .INP(n39), .Z(n6804) );
  NBUFFX2 U1743 ( .INP(n38), .Z(n6793) );
  NBUFFX2 U1744 ( .INP(n37), .Z(n6782) );
  NBUFFX2 U1745 ( .INP(n36), .Z(n6771) );
  NBUFFX2 U1746 ( .INP(n35), .Z(n6760) );
  NBUFFX2 U1747 ( .INP(n34), .Z(n6749) );
  NBUFFX2 U1748 ( .INP(n41), .Z(n6825) );
  NBUFFX2 U1749 ( .INP(n40), .Z(n6814) );
  NBUFFX2 U1750 ( .INP(n39), .Z(n6803) );
  NBUFFX2 U1751 ( .INP(n38), .Z(n6792) );
  NBUFFX2 U1752 ( .INP(n37), .Z(n6781) );
  NBUFFX2 U1753 ( .INP(n36), .Z(n6770) );
  NBUFFX2 U1754 ( .INP(n35), .Z(n6759) );
  NBUFFX2 U1755 ( .INP(n34), .Z(n6748) );
  NBUFFX2 U1756 ( .INP(n41), .Z(n6824) );
  NBUFFX2 U1757 ( .INP(n40), .Z(n6813) );
  NBUFFX2 U1758 ( .INP(n39), .Z(n6802) );
  NBUFFX2 U1759 ( .INP(n38), .Z(n6791) );
  NBUFFX2 U1769 ( .INP(n37), .Z(n6780) );
  NBUFFX2 U1770 ( .INP(n36), .Z(n6769) );
  NBUFFX2 U1771 ( .INP(n35), .Z(n6758) );
  NBUFFX2 U1772 ( .INP(n34), .Z(n6747) );
  NBUFFX2 U1773 ( .INP(n41), .Z(n6823) );
  NBUFFX2 U1774 ( .INP(n40), .Z(n6812) );
  NBUFFX2 U1775 ( .INP(n39), .Z(n6801) );
  NBUFFX2 U1776 ( .INP(n38), .Z(n6790) );
  NBUFFX2 U1777 ( .INP(n37), .Z(n6779) );
  NBUFFX2 U1778 ( .INP(n36), .Z(n6768) );
  NBUFFX2 U1779 ( .INP(n35), .Z(n6757) );
  NBUFFX2 U1780 ( .INP(n34), .Z(n6746) );
  NBUFFX2 U1781 ( .INP(n41), .Z(n6822) );
  NBUFFX2 U1782 ( .INP(n40), .Z(n6811) );
  NBUFFX2 U1783 ( .INP(n39), .Z(n6800) );
  NBUFFX2 U1784 ( .INP(n38), .Z(n6789) );
  NBUFFX2 U1785 ( .INP(n37), .Z(n6778) );
  NBUFFX2 U1786 ( .INP(n36), .Z(n6767) );
  NBUFFX2 U1787 ( .INP(n35), .Z(n6756) );
  NBUFFX2 U1788 ( .INP(n34), .Z(n6745) );
  NBUFFX2 U1789 ( .INP(n41), .Z(n6821) );
  NBUFFX2 U1790 ( .INP(n40), .Z(n6810) );
  NBUFFX2 U1791 ( .INP(n39), .Z(n6799) );
  NBUFFX2 U1792 ( .INP(n38), .Z(n6788) );
  NBUFFX2 U1868 ( .INP(n37), .Z(n6777) );
  NBUFFX2 U1869 ( .INP(n36), .Z(n6766) );
  NBUFFX2 U1870 ( .INP(n35), .Z(n6755) );
  NBUFFX2 U1871 ( .INP(n34), .Z(n6744) );
  NBUFFX2 U1872 ( .INP(n41), .Z(n6820) );
  NBUFFX2 U1873 ( .INP(n40), .Z(n6809) );
  NBUFFX2 U1874 ( .INP(n39), .Z(n6798) );
  NBUFFX2 U1875 ( .INP(n38), .Z(n6787) );
  NBUFFX2 U1876 ( .INP(n37), .Z(n6776) );
  NBUFFX2 U1877 ( .INP(n36), .Z(n6765) );
  NBUFFX2 U1878 ( .INP(n35), .Z(n6754) );
  NBUFFX2 U1879 ( .INP(n34), .Z(n6743) );
  NBUFFX2 U1880 ( .INP(n41), .Z(n6819) );
  NBUFFX2 U1881 ( .INP(n40), .Z(n6808) );
  NBUFFX2 U1882 ( .INP(n39), .Z(n6797) );
  NBUFFX2 U1883 ( .INP(n38), .Z(n6786) );
  NBUFFX2 U1884 ( .INP(n37), .Z(n6775) );
  NBUFFX2 U1885 ( .INP(n36), .Z(n6764) );
  NBUFFX2 U1886 ( .INP(n35), .Z(n6753) );
  NBUFFX2 U1887 ( .INP(n34), .Z(n6742) );
  NBUFFX2 U1888 ( .INP(n41), .Z(n6818) );
  NBUFFX2 U1889 ( .INP(n40), .Z(n6807) );
  NBUFFX2 U1890 ( .INP(n39), .Z(n6796) );
  NBUFFX2 U1891 ( .INP(n38), .Z(n6785) );
  NBUFFX2 U1892 ( .INP(n37), .Z(n6774) );
  NBUFFX2 U1902 ( .INP(n36), .Z(n6763) );
  NBUFFX2 U1903 ( .INP(n35), .Z(n6752) );
  NBUFFX2 U1904 ( .INP(n34), .Z(n6741) );
  NBUFFX2 U1905 ( .INP(n50), .Z(n7004) );
  NBUFFX2 U1906 ( .INP(n27), .Z(n6993) );
  NBUFFX2 U1907 ( .INP(n26), .Z(n6982) );
  NBUFFX2 U1908 ( .INP(n25), .Z(n6971) );
  NBUFFX2 U1909 ( .INP(n24), .Z(n6894) );
  NBUFFX2 U1910 ( .INP(n23), .Z(n6883) );
  NBUFFX2 U1911 ( .INP(n51), .Z(n6872) );
  NBUFFX2 U1912 ( .INP(n22), .Z(n6861) );
  NBUFFX2 U1913 ( .INP(n21), .Z(n6850) );
  NBUFFX2 U1914 ( .INP(n20), .Z(n6839) );
  NBUFFX2 U1915 ( .INP(n33), .Z(n6960) );
  NBUFFX2 U1916 ( .INP(n32), .Z(n6949) );
  NBUFFX2 U1917 ( .INP(n31), .Z(n6938) );
  NBUFFX2 U1918 ( .INP(n30), .Z(n6927) );
  NBUFFX2 U1919 ( .INP(n29), .Z(n6916) );
  NBUFFX2 U1920 ( .INP(n28), .Z(n6905) );
  NBUFFX2 U1921 ( .INP(n41), .Z(n6828) );
  NBUFFX2 U1922 ( .INP(n40), .Z(n6817) );
  NBUFFX2 U1923 ( .INP(n39), .Z(n6806) );
  NBUFFX2 U1924 ( .INP(n38), .Z(n6795) );
  NBUFFX2 U1925 ( .INP(n37), .Z(n6784) );
  NBUFFX2 U1942 ( .INP(n36), .Z(n6773) );
  NBUFFX2 U1954 ( .INP(n35), .Z(n6762) );
  NBUFFX2 U1976 ( .INP(n34), .Z(n6751) );
  NBUFFX2 U1989 ( .INP(n49), .Z(n7098) );
  NBUFFX2 U2001 ( .INP(n48), .Z(n7081) );
  NBUFFX2 U2002 ( .INP(n47), .Z(n7070) );
  NBUFFX2 U2003 ( .INP(n46), .Z(n7059) );
  NBUFFX2 U2004 ( .INP(n45), .Z(n7048) );
  NBUFFX2 U2005 ( .INP(n44), .Z(n7037) );
  NBUFFX2 U2006 ( .INP(n43), .Z(n7026) );
  NBUFFX2 U2007 ( .INP(n42), .Z(n7015) );
  NBUFFX2 U2008 ( .INP(n5969), .Z(n5896) );
  NBUFFX2 U2009 ( .INP(n5972), .Z(n5895) );
  NBUFFX2 U2010 ( .INP(n5972), .Z(n5894) );
  NBUFFX2 U2011 ( .INP(n5972), .Z(n5893) );
  NBUFFX2 U2012 ( .INP(n5971), .Z(n5892) );
  NBUFFX2 U2013 ( .INP(n5971), .Z(n5891) );
  NBUFFX2 U2014 ( .INP(n5971), .Z(n5890) );
  NBUFFX2 U2015 ( .INP(n5970), .Z(n5889) );
  NBUFFX2 U2016 ( .INP(n5970), .Z(n5888) );
  NBUFFX2 U2017 ( .INP(n5970), .Z(n5887) );
  NBUFFX2 U2018 ( .INP(n5969), .Z(n5886) );
  NBUFFX2 U2019 ( .INP(n5969), .Z(n5885) );
  NBUFFX2 U2020 ( .INP(n5969), .Z(n5884) );
  NBUFFX2 U2021 ( .INP(n5968), .Z(n5883) );
  NBUFFX2 U2022 ( .INP(n5968), .Z(n5882) );
  NBUFFX2 U2023 ( .INP(n5968), .Z(n5881) );
  NBUFFX2 U2024 ( .INP(n5967), .Z(n5880) );
  NBUFFX2 U2034 ( .INP(n5967), .Z(n5879) );
  NBUFFX2 U2035 ( .INP(n5967), .Z(n5878) );
  NBUFFX2 U2036 ( .INP(n5966), .Z(n5877) );
  NBUFFX2 U2037 ( .INP(n5966), .Z(n5876) );
  NBUFFX2 U2038 ( .INP(n5966), .Z(n5875) );
  NBUFFX2 U2039 ( .INP(n5965), .Z(n5874) );
  NBUFFX2 U2040 ( .INP(n5788), .Z(n5790) );
  NBUFFX2 U2041 ( .INP(n5788), .Z(n5791) );
  NBUFFX2 U2042 ( .INP(n5787), .Z(n5800) );
  NBUFFX2 U2043 ( .INP(n5787), .Z(n5801) );
  NBUFFX2 U2044 ( .INP(n5786), .Z(n5812) );
  NBUFFX2 U2045 ( .INP(n5786), .Z(n5813) );
  NBUFFX2 U2046 ( .INP(n5785), .Z(n5824) );
  NBUFFX2 U2047 ( .INP(n5785), .Z(n5825) );
  NBUFFX2 U2048 ( .INP(n5784), .Z(n5836) );
  NBUFFX2 U2049 ( .INP(n5784), .Z(n5837) );
  NBUFFX2 U2050 ( .INP(n5783), .Z(n5848) );
  NBUFFX2 U2051 ( .INP(n5783), .Z(n5849) );
  NBUFFX2 U2052 ( .INP(n5782), .Z(n5860) );
  NBUFFX2 U2053 ( .INP(n5782), .Z(n5861) );
  NBUFFX2 U2054 ( .INP(n5788), .Z(n5792) );
  NBUFFX2 U2055 ( .INP(n5788), .Z(n5793) );
  NBUFFX2 U2056 ( .INP(n5788), .Z(n5794) );
  NBUFFX2 U2057 ( .INP(n5788), .Z(n5795) );
  NBUFFX2 U2109 ( .INP(n5788), .Z(n5796) );
  NBUFFX2 U2122 ( .INP(n5788), .Z(n5797) );
  NBUFFX2 U2133 ( .INP(n5788), .Z(n5798) );
  NBUFFX2 U2134 ( .INP(n5788), .Z(n5799) );
  NBUFFX2 U2135 ( .INP(n5787), .Z(n5802) );
  NBUFFX2 U2136 ( .INP(n5787), .Z(n5803) );
  NBUFFX2 U2137 ( .INP(n5787), .Z(n5804) );
  NBUFFX2 U2138 ( .INP(n5787), .Z(n5805) );
  NBUFFX2 U2139 ( .INP(n5787), .Z(n5806) );
  NBUFFX2 U2140 ( .INP(n5787), .Z(n5807) );
  NBUFFX2 U2141 ( .INP(n5787), .Z(n5808) );
  NBUFFX2 U2142 ( .INP(n5787), .Z(n5809) );
  NBUFFX2 U2143 ( .INP(n5787), .Z(n5810) );
  NBUFFX2 U2144 ( .INP(n5787), .Z(n5811) );
  NBUFFX2 U2145 ( .INP(n5786), .Z(n5814) );
  NBUFFX2 U2146 ( .INP(n5786), .Z(n5815) );
  NBUFFX2 U2147 ( .INP(n5786), .Z(n5816) );
  NBUFFX2 U2148 ( .INP(n5786), .Z(n5817) );
  NBUFFX2 U2149 ( .INP(n5786), .Z(n5818) );
  NBUFFX2 U2150 ( .INP(n5786), .Z(n5819) );
  NBUFFX2 U2151 ( .INP(n5786), .Z(n5820) );
  NBUFFX2 U2152 ( .INP(n5786), .Z(n5821) );
  NBUFFX2 U2153 ( .INP(n5786), .Z(n5822) );
  NBUFFX2 U2154 ( .INP(n5786), .Z(n5823) );
  NBUFFX2 U2155 ( .INP(n5785), .Z(n5826) );
  NBUFFX2 U2156 ( .INP(n5785), .Z(n5827) );
  NBUFFX2 U2166 ( .INP(n5785), .Z(n5828) );
  NBUFFX2 U2167 ( .INP(n5785), .Z(n5829) );
  NBUFFX2 U2168 ( .INP(n5785), .Z(n5830) );
  NBUFFX2 U2169 ( .INP(n5785), .Z(n5831) );
  NBUFFX2 U2170 ( .INP(n5785), .Z(n5832) );
  NBUFFX2 U2171 ( .INP(n5785), .Z(n5833) );
  NBUFFX2 U2172 ( .INP(n5785), .Z(n5834) );
  NBUFFX2 U2173 ( .INP(n5785), .Z(n5835) );
  NBUFFX2 U2174 ( .INP(n5784), .Z(n5838) );
  NBUFFX2 U2175 ( .INP(n5784), .Z(n5839) );
  NBUFFX2 U2176 ( .INP(n5784), .Z(n5840) );
  NBUFFX2 U2177 ( .INP(n5784), .Z(n5841) );
  NBUFFX2 U2178 ( .INP(n5784), .Z(n5842) );
  NBUFFX2 U2179 ( .INP(n5784), .Z(n5843) );
  NBUFFX2 U2180 ( .INP(n5784), .Z(n5844) );
  NBUFFX2 U2181 ( .INP(n5784), .Z(n5845) );
  NBUFFX2 U2182 ( .INP(n5784), .Z(n5846) );
  NBUFFX2 U2183 ( .INP(n5784), .Z(n5847) );
  NBUFFX2 U2184 ( .INP(n5783), .Z(n5850) );
  NBUFFX2 U2185 ( .INP(n5783), .Z(n5851) );
  NBUFFX2 U2186 ( .INP(n5783), .Z(n5852) );
  NBUFFX2 U2187 ( .INP(n5783), .Z(n5853) );
  NBUFFX2 U2188 ( .INP(n5783), .Z(n5854) );
  NBUFFX2 U2189 ( .INP(n5783), .Z(n5855) );
  NBUFFX2 U2265 ( .INP(n5783), .Z(n5856) );
  NBUFFX2 U2266 ( .INP(n5783), .Z(n5857) );
  NBUFFX2 U2267 ( .INP(n5783), .Z(n5858) );
  NBUFFX2 U2268 ( .INP(n5783), .Z(n5859) );
  NBUFFX2 U2269 ( .INP(n5782), .Z(n5862) );
  NBUFFX2 U2270 ( .INP(n5782), .Z(n5863) );
  NBUFFX2 U2271 ( .INP(n5782), .Z(n5864) );
  NBUFFX2 U2272 ( .INP(n5782), .Z(n5865) );
  NBUFFX2 U2273 ( .INP(n5782), .Z(n5866) );
  NBUFFX2 U2274 ( .INP(n5782), .Z(n5867) );
  NBUFFX2 U2275 ( .INP(n5782), .Z(n5868) );
  NBUFFX2 U2276 ( .INP(n5782), .Z(n5869) );
  NBUFFX2 U2277 ( .INP(n5782), .Z(n5870) );
  NBUFFX2 U2278 ( .INP(n5782), .Z(n5871) );
  NBUFFX2 U2279 ( .INP(n5788), .Z(n5872) );
  NBUFFX2 U2280 ( .INP(n5785), .Z(n5873) );
  NBUFFX2 U2281 ( .INP(n5756), .Z(n5736) );
  NBUFFX2 U2282 ( .INP(n5756), .Z(n5737) );
  NBUFFX2 U2283 ( .INP(n5756), .Z(n5738) );
  NBUFFX2 U2284 ( .INP(n5756), .Z(n5739) );
  NBUFFX2 U2285 ( .INP(n5757), .Z(n5744) );
  NBUFFX2 U2286 ( .INP(n5757), .Z(n5745) );
  INVX0 U2287 ( .INP(n204), .ZN(n7103) );
  INVX0 U2288 ( .INP(n204), .ZN(n7102) );
  INVX0 U2298 ( .INP(n204), .ZN(n7101) );
  NBUFFX2 U2299 ( .INP(n5756), .Z(n5740) );
  NBUFFX2 U2300 ( .INP(n5756), .Z(n5741) );
  NBUFFX2 U2301 ( .INP(n5756), .Z(n5742) );
  NBUFFX2 U2302 ( .INP(n5756), .Z(n5743) );
  NBUFFX2 U2303 ( .INP(n5757), .Z(n5746) );
  NBUFFX2 U2304 ( .INP(n5757), .Z(n5747) );
  NBUFFX2 U2305 ( .INP(n5757), .Z(n5748) );
  NBUFFX2 U2306 ( .INP(n5757), .Z(n5749) );
  NBUFFX2 U2307 ( .INP(n5757), .Z(n5750) );
  NBUFFX2 U2308 ( .INP(n5757), .Z(n5751) );
  NBUFFX2 U2309 ( .INP(n5757), .Z(n5752) );
  NBUFFX2 U2310 ( .INP(n5757), .Z(n5753) );
  NBUFFX2 U2311 ( .INP(n5757), .Z(n5754) );
  NBUFFX2 U2312 ( .INP(n5757), .Z(n5755) );
  NBUFFX2 U2313 ( .INP(n5788), .Z(n5789) );
  NBUFFX2 U2314 ( .INP(n5756), .Z(n5735) );
  NBUFFX2 U2315 ( .INP(n7359), .Z(n5974) );
  NBUFFX2 U2316 ( .INP(n7359), .Z(n5975) );
  NBUFFX2 U2317 ( .INP(n7359), .Z(n5973) );
  NBUFFX2 U2318 ( .INP(n7356), .Z(n7357) );
  NBUFFX2 U2319 ( .INP(n7355), .Z(n7356) );
  NBUFFX2 U2320 ( .INP(n7354), .Z(n7355) );
  NBUFFX2 U2321 ( .INP(n7358), .Z(n7354) );
  NBUFFX2 U2397 ( .INP(n7358), .Z(n7353) );
  AND4X1 U2398 ( .IN1(wraddr[6]), .IN2(n270), .IN3(n7366), .IN4(n7367), .Q(
        n306) );
  AND4X1 U2399 ( .IN1(wraddr[4]), .IN2(n270), .IN3(n7367), .IN4(n7368), .Q(
        n357) );
  NOR2X0 U2400 ( .IN1(n7363), .IN2(wraddr[0]), .QN(n378) );
  NOR2X0 U2401 ( .IN1(n7365), .IN2(wraddr[2]), .QN(n384) );
  INVX0 U2402 ( .INP(wraddr[4]), .ZN(n7366) );
  AO22X1 U2403 ( .IN1(n7097), .IN2(n6647), .IN3(\FIFO[111][0] ), .IN4(n6648), 
        .Q(n979) );
  AO22X1 U2404 ( .IN1(n7080), .IN2(n6647), .IN3(\FIFO[111][1] ), .IN4(n6648), 
        .Q(n980) );
  AO22X1 U2405 ( .IN1(n7069), .IN2(n6647), .IN3(\FIFO[111][2] ), .IN4(n6648), 
        .Q(n981) );
  AO22X1 U2406 ( .IN1(n7058), .IN2(n6647), .IN3(\FIFO[111][3] ), .IN4(n6648), 
        .Q(n982) );
  AO22X1 U2407 ( .IN1(n7047), .IN2(n6647), .IN3(\FIFO[111][4] ), .IN4(n6648), 
        .Q(n983) );
  AO22X1 U2408 ( .IN1(n7036), .IN2(n6647), .IN3(\FIFO[111][5] ), .IN4(n6648), 
        .Q(n984) );
  AO22X1 U2409 ( .IN1(n7025), .IN2(n6647), .IN3(\FIFO[111][6] ), .IN4(n6648), 
        .Q(n985) );
  AO22X1 U2410 ( .IN1(n7014), .IN2(n6646), .IN3(\FIFO[111][7] ), .IN4(n6648), 
        .Q(n986) );
  AO22X1 U2411 ( .IN1(n7003), .IN2(n6646), .IN3(\FIFO[111][8] ), .IN4(n6648), 
        .Q(n987) );
  AO22X1 U2412 ( .IN1(n6992), .IN2(n6646), .IN3(\FIFO[111][9] ), .IN4(n6648), 
        .Q(n988) );
  AO22X1 U2413 ( .IN1(n6981), .IN2(n6646), .IN3(\FIFO[111][10] ), .IN4(n6648), 
        .Q(n989) );
  AO22X1 U2414 ( .IN1(n6970), .IN2(n6646), .IN3(\FIFO[111][11] ), .IN4(n6648), 
        .Q(n990) );
  AO22X1 U2415 ( .IN1(n6959), .IN2(n6646), .IN3(\FIFO[111][12] ), .IN4(n6649), 
        .Q(n991) );
  AO22X1 U2416 ( .IN1(n6948), .IN2(n6646), .IN3(\FIFO[111][13] ), .IN4(n6649), 
        .Q(n992) );
  AO22X1 U2417 ( .IN1(n6937), .IN2(n6645), .IN3(\FIFO[111][14] ), .IN4(n6649), 
        .Q(n993) );
  AO22X1 U2418 ( .IN1(n6926), .IN2(n6645), .IN3(\FIFO[111][15] ), .IN4(n6649), 
        .Q(n994) );
  AO22X1 U2419 ( .IN1(n6915), .IN2(n6645), .IN3(\FIFO[111][16] ), .IN4(n6649), 
        .Q(n995) );
  AO22X1 U2420 ( .IN1(n6904), .IN2(n6645), .IN3(\FIFO[111][17] ), .IN4(n6649), 
        .Q(n996) );
  AO22X1 U2421 ( .IN1(n6893), .IN2(n6645), .IN3(\FIFO[111][18] ), .IN4(n6649), 
        .Q(n997) );
  AO22X1 U2431 ( .IN1(n6882), .IN2(n6645), .IN3(\FIFO[111][19] ), .IN4(n6649), 
        .Q(n998) );
  AO22X1 U2432 ( .IN1(n6871), .IN2(n6645), .IN3(\FIFO[111][20] ), .IN4(n6649), 
        .Q(n999) );
  AO22X1 U2433 ( .IN1(n6860), .IN2(n6647), .IN3(\FIFO[111][21] ), .IN4(n6649), 
        .Q(n1000) );
  AO22X1 U2434 ( .IN1(n6849), .IN2(n6646), .IN3(\FIFO[111][22] ), .IN4(n6649), 
        .Q(n1001) );
  AO22X1 U2435 ( .IN1(n6838), .IN2(n6645), .IN3(\FIFO[111][23] ), .IN4(n6649), 
        .Q(n1002) );
  AO22X1 U2436 ( .IN1(n7097), .IN2(n6641), .IN3(\FIFO[110][0] ), .IN4(n6642), 
        .Q(n1011) );
  AO22X1 U2437 ( .IN1(n7080), .IN2(n6641), .IN3(\FIFO[110][1] ), .IN4(n6642), 
        .Q(n1012) );
  AO22X1 U2438 ( .IN1(n7069), .IN2(n6641), .IN3(\FIFO[110][2] ), .IN4(n6642), 
        .Q(n1013) );
  AO22X1 U2439 ( .IN1(n7058), .IN2(n6641), .IN3(\FIFO[110][3] ), .IN4(n6642), 
        .Q(n1014) );
  AO22X1 U2440 ( .IN1(n7047), .IN2(n6641), .IN3(\FIFO[110][4] ), .IN4(n6642), 
        .Q(n1015) );
  AO22X1 U2441 ( .IN1(n7036), .IN2(n6641), .IN3(\FIFO[110][5] ), .IN4(n6642), 
        .Q(n1016) );
  AO22X1 U2442 ( .IN1(n7025), .IN2(n6641), .IN3(\FIFO[110][6] ), .IN4(n6642), 
        .Q(n1017) );
  AO22X1 U2443 ( .IN1(n7014), .IN2(n6640), .IN3(\FIFO[110][7] ), .IN4(n6642), 
        .Q(n1018) );
  AO22X1 U2444 ( .IN1(n7003), .IN2(n6640), .IN3(\FIFO[110][8] ), .IN4(n6642), 
        .Q(n1019) );
  AO22X1 U2445 ( .IN1(n6992), .IN2(n6640), .IN3(\FIFO[110][9] ), .IN4(n6642), 
        .Q(n1020) );
  AO22X1 U2446 ( .IN1(n6981), .IN2(n6640), .IN3(\FIFO[110][10] ), .IN4(n6642), 
        .Q(n1021) );
  AO22X1 U2447 ( .IN1(n6970), .IN2(n6640), .IN3(\FIFO[110][11] ), .IN4(n6642), 
        .Q(n1022) );
  AO22X1 U2448 ( .IN1(n6959), .IN2(n6640), .IN3(\FIFO[110][12] ), .IN4(n6643), 
        .Q(n1023) );
  AO22X1 U2449 ( .IN1(n6948), .IN2(n6640), .IN3(\FIFO[110][13] ), .IN4(n6643), 
        .Q(n1024) );
  AO22X1 U2450 ( .IN1(n6937), .IN2(n6639), .IN3(\FIFO[110][14] ), .IN4(n6643), 
        .Q(n1025) );
  AO22X1 U2451 ( .IN1(n6926), .IN2(n6639), .IN3(\FIFO[110][15] ), .IN4(n6643), 
        .Q(n1026) );
  AO22X1 U2452 ( .IN1(n6915), .IN2(n6639), .IN3(\FIFO[110][16] ), .IN4(n6643), 
        .Q(n1027) );
  AO22X1 U2453 ( .IN1(n6904), .IN2(n6639), .IN3(\FIFO[110][17] ), .IN4(n6643), 
        .Q(n1028) );
  AO22X1 U2454 ( .IN1(n6893), .IN2(n6639), .IN3(\FIFO[110][18] ), .IN4(n6643), 
        .Q(n1029) );
  AO22X1 U2496 ( .IN1(n6882), .IN2(n6639), .IN3(\FIFO[110][19] ), .IN4(n6643), 
        .Q(n1030) );
  AO22X1 U2530 ( .IN1(n6871), .IN2(n6639), .IN3(\FIFO[110][20] ), .IN4(n6643), 
        .Q(n1031) );
  AO22X1 U2531 ( .IN1(n6860), .IN2(n6641), .IN3(\FIFO[110][21] ), .IN4(n6643), 
        .Q(n1032) );
  AO22X1 U2532 ( .IN1(n6849), .IN2(n6640), .IN3(\FIFO[110][22] ), .IN4(n6643), 
        .Q(n1033) );
  AO22X1 U2533 ( .IN1(n6838), .IN2(n6639), .IN3(\FIFO[110][23] ), .IN4(n6643), 
        .Q(n1034) );
  AO22X1 U2534 ( .IN1(n7096), .IN2(n6623), .IN3(\FIFO[107][0] ), .IN4(n6624), 
        .Q(n1107) );
  AO22X1 U2535 ( .IN1(n7079), .IN2(n6622), .IN3(\FIFO[107][1] ), .IN4(n6624), 
        .Q(n1108) );
  AO22X1 U2536 ( .IN1(n7068), .IN2(n6621), .IN3(\FIFO[107][2] ), .IN4(n6624), 
        .Q(n1109) );
  AO22X1 U2537 ( .IN1(n7057), .IN2(n6623), .IN3(\FIFO[107][3] ), .IN4(n6624), 
        .Q(n1110) );
  AO22X1 U2538 ( .IN1(n7046), .IN2(n6622), .IN3(\FIFO[107][4] ), .IN4(n6624), 
        .Q(n1111) );
  AO22X1 U2539 ( .IN1(n7035), .IN2(n6621), .IN3(\FIFO[107][5] ), .IN4(n6624), 
        .Q(n1112) );
  AO22X1 U2540 ( .IN1(n7024), .IN2(n6623), .IN3(\FIFO[107][6] ), .IN4(n6624), 
        .Q(n1113) );
  AO22X1 U2541 ( .IN1(n7013), .IN2(n6623), .IN3(\FIFO[107][7] ), .IN4(n6624), 
        .Q(n1114) );
  AO22X1 U2542 ( .IN1(n7002), .IN2(n6623), .IN3(\FIFO[107][8] ), .IN4(n6624), 
        .Q(n1115) );
  AO22X1 U2543 ( .IN1(n6991), .IN2(n6623), .IN3(\FIFO[107][9] ), .IN4(n6624), 
        .Q(n1116) );
  AO22X1 U2544 ( .IN1(n6980), .IN2(n6623), .IN3(\FIFO[107][10] ), .IN4(n6624), 
        .Q(n1117) );
  AO22X1 U2545 ( .IN1(n6969), .IN2(n6623), .IN3(\FIFO[107][11] ), .IN4(n6624), 
        .Q(n1118) );
  AO22X1 U2546 ( .IN1(n6958), .IN2(n6623), .IN3(\FIFO[107][12] ), .IN4(n6625), 
        .Q(n1119) );
  AO22X1 U2547 ( .IN1(n6947), .IN2(n6623), .IN3(\FIFO[107][13] ), .IN4(n6625), 
        .Q(n1120) );
  AO22X1 U2548 ( .IN1(n6936), .IN2(n6622), .IN3(\FIFO[107][14] ), .IN4(n6625), 
        .Q(n1121) );
  AO22X1 U2549 ( .IN1(n6925), .IN2(n6622), .IN3(\FIFO[107][15] ), .IN4(n6625), 
        .Q(n1122) );
  AO22X1 U2550 ( .IN1(n6914), .IN2(n6622), .IN3(\FIFO[107][16] ), .IN4(n6625), 
        .Q(n1123) );
  AO22X1 U2551 ( .IN1(n6903), .IN2(n6622), .IN3(\FIFO[107][17] ), .IN4(n6625), 
        .Q(n1124) );
  AO22X1 U2552 ( .IN1(n6892), .IN2(n6622), .IN3(\FIFO[107][18] ), .IN4(n6625), 
        .Q(n1125) );
  AO22X1 U2553 ( .IN1(n6881), .IN2(n6622), .IN3(\FIFO[107][19] ), .IN4(n6625), 
        .Q(n1126) );
  AO22X1 U2563 ( .IN1(n6870), .IN2(n6622), .IN3(\FIFO[107][20] ), .IN4(n6625), 
        .Q(n1127) );
  AO22X1 U2564 ( .IN1(n6859), .IN2(n6621), .IN3(\FIFO[107][21] ), .IN4(n6625), 
        .Q(n1128) );
  AO22X1 U2565 ( .IN1(n6848), .IN2(n6621), .IN3(\FIFO[107][22] ), .IN4(n6625), 
        .Q(n1129) );
  AO22X1 U2566 ( .IN1(n6837), .IN2(n6621), .IN3(\FIFO[107][23] ), .IN4(n6625), 
        .Q(n1130) );
  AO22X1 U2567 ( .IN1(n7096), .IN2(n6617), .IN3(\FIFO[106][0] ), .IN4(n6618), 
        .Q(n1139) );
  AO22X1 U2568 ( .IN1(n7079), .IN2(n6617), .IN3(\FIFO[106][1] ), .IN4(n6618), 
        .Q(n1140) );
  AO22X1 U2569 ( .IN1(n7068), .IN2(n6617), .IN3(\FIFO[106][2] ), .IN4(n6618), 
        .Q(n1141) );
  AO22X1 U2570 ( .IN1(n7057), .IN2(n6617), .IN3(\FIFO[106][3] ), .IN4(n6618), 
        .Q(n1142) );
  AO22X1 U2571 ( .IN1(n7046), .IN2(n6617), .IN3(\FIFO[106][4] ), .IN4(n6618), 
        .Q(n1143) );
  AO22X1 U2572 ( .IN1(n7035), .IN2(n6617), .IN3(\FIFO[106][5] ), .IN4(n6618), 
        .Q(n1144) );
  AO22X1 U2573 ( .IN1(n7024), .IN2(n6617), .IN3(\FIFO[106][6] ), .IN4(n6618), 
        .Q(n1145) );
  AO22X1 U2574 ( .IN1(n7013), .IN2(n6616), .IN3(\FIFO[106][7] ), .IN4(n6618), 
        .Q(n1146) );
  AO22X1 U2575 ( .IN1(n7002), .IN2(n6616), .IN3(\FIFO[106][8] ), .IN4(n6618), 
        .Q(n1147) );
  AO22X1 U2576 ( .IN1(n6991), .IN2(n6616), .IN3(\FIFO[106][9] ), .IN4(n6618), 
        .Q(n1148) );
  AO22X1 U2577 ( .IN1(n6980), .IN2(n6616), .IN3(\FIFO[106][10] ), .IN4(n6618), 
        .Q(n1149) );
  AO22X1 U2578 ( .IN1(n6969), .IN2(n6616), .IN3(\FIFO[106][11] ), .IN4(n6618), 
        .Q(n1150) );
  AO22X1 U2579 ( .IN1(n6958), .IN2(n6616), .IN3(\FIFO[106][12] ), .IN4(n6619), 
        .Q(n1151) );
  AO22X1 U2580 ( .IN1(n6947), .IN2(n6616), .IN3(\FIFO[106][13] ), .IN4(n6619), 
        .Q(n1152) );
  AO22X1 U2581 ( .IN1(n6936), .IN2(n6615), .IN3(\FIFO[106][14] ), .IN4(n6619), 
        .Q(n1153) );
  AO22X1 U2582 ( .IN1(n6925), .IN2(n6615), .IN3(\FIFO[106][15] ), .IN4(n6619), 
        .Q(n1154) );
  AO22X1 U2583 ( .IN1(n6914), .IN2(n6615), .IN3(\FIFO[106][16] ), .IN4(n6619), 
        .Q(n1155) );
  AO22X1 U2584 ( .IN1(n6903), .IN2(n6615), .IN3(\FIFO[106][17] ), .IN4(n6619), 
        .Q(n1156) );
  AO22X1 U2585 ( .IN1(n6892), .IN2(n6615), .IN3(\FIFO[106][18] ), .IN4(n6619), 
        .Q(n1157) );
  AO22X1 U2586 ( .IN1(n6881), .IN2(n6615), .IN3(\FIFO[106][19] ), .IN4(n6619), 
        .Q(n1158) );
  AO22X1 U2598 ( .IN1(n6870), .IN2(n6615), .IN3(\FIFO[106][20] ), .IN4(n6619), 
        .Q(n1159) );
  AO22X1 U2613 ( .IN1(n6859), .IN2(n6617), .IN3(\FIFO[106][21] ), .IN4(n6619), 
        .Q(n1160) );
  AO22X1 U2662 ( .IN1(n6848), .IN2(n6616), .IN3(\FIFO[106][22] ), .IN4(n6619), 
        .Q(n1161) );
  AO22X1 U2663 ( .IN1(n6837), .IN2(n6615), .IN3(\FIFO[106][23] ), .IN4(n6619), 
        .Q(n1162) );
  AO22X1 U2664 ( .IN1(n7096), .IN2(n6599), .IN3(\FIFO[103][0] ), .IN4(n6600), 
        .Q(n1235) );
  AO22X1 U2665 ( .IN1(n7079), .IN2(n6599), .IN3(\FIFO[103][1] ), .IN4(n6600), 
        .Q(n1236) );
  AO22X1 U2666 ( .IN1(n7068), .IN2(n6599), .IN3(\FIFO[103][2] ), .IN4(n6600), 
        .Q(n1237) );
  AO22X1 U2667 ( .IN1(n7057), .IN2(n6599), .IN3(\FIFO[103][3] ), .IN4(n6600), 
        .Q(n1238) );
  AO22X1 U2668 ( .IN1(n7046), .IN2(n6599), .IN3(\FIFO[103][4] ), .IN4(n6600), 
        .Q(n1239) );
  AO22X1 U2669 ( .IN1(n7035), .IN2(n6599), .IN3(\FIFO[103][5] ), .IN4(n6600), 
        .Q(n1240) );
  AO22X1 U2670 ( .IN1(n7024), .IN2(n6599), .IN3(\FIFO[103][6] ), .IN4(n6600), 
        .Q(n1241) );
  AO22X1 U2671 ( .IN1(n7013), .IN2(n6598), .IN3(\FIFO[103][7] ), .IN4(n6600), 
        .Q(n1242) );
  AO22X1 U2672 ( .IN1(n7002), .IN2(n6598), .IN3(\FIFO[103][8] ), .IN4(n6600), 
        .Q(n1243) );
  AO22X1 U2673 ( .IN1(n6991), .IN2(n6598), .IN3(\FIFO[103][9] ), .IN4(n6600), 
        .Q(n1244) );
  AO22X1 U2674 ( .IN1(n6980), .IN2(n6598), .IN3(\FIFO[103][10] ), .IN4(n6600), 
        .Q(n1245) );
  AO22X1 U2675 ( .IN1(n6969), .IN2(n6598), .IN3(\FIFO[103][11] ), .IN4(n6600), 
        .Q(n1246) );
  AO22X1 U2676 ( .IN1(n6947), .IN2(n6598), .IN3(\FIFO[103][13] ), .IN4(n6601), 
        .Q(n1248) );
  AO22X1 U2677 ( .IN1(n6936), .IN2(n6599), .IN3(\FIFO[103][14] ), .IN4(n6601), 
        .Q(n1249) );
  AO22X1 U2678 ( .IN1(n6925), .IN2(n6598), .IN3(\FIFO[103][15] ), .IN4(n6601), 
        .Q(n1250) );
  AO22X1 U2679 ( .IN1(n6914), .IN2(n6597), .IN3(\FIFO[103][16] ), .IN4(n6601), 
        .Q(n1251) );
  AO22X1 U2680 ( .IN1(n6903), .IN2(n6599), .IN3(\FIFO[103][17] ), .IN4(n6601), 
        .Q(n1252) );
  AO22X1 U2681 ( .IN1(n6892), .IN2(n6598), .IN3(\FIFO[103][18] ), .IN4(n6601), 
        .Q(n1253) );
  AO22X1 U2682 ( .IN1(n6881), .IN2(n6597), .IN3(\FIFO[103][19] ), .IN4(n6601), 
        .Q(n1254) );
  AO22X1 U2683 ( .IN1(n6870), .IN2(n6599), .IN3(\FIFO[103][20] ), .IN4(n6601), 
        .Q(n1255) );
  AO22X1 U2684 ( .IN1(n6859), .IN2(n6597), .IN3(\FIFO[103][21] ), .IN4(n6601), 
        .Q(n1256) );
  AO22X1 U2685 ( .IN1(n6848), .IN2(n6597), .IN3(\FIFO[103][22] ), .IN4(n6601), 
        .Q(n1257) );
  AO22X1 U2695 ( .IN1(n6837), .IN2(n6597), .IN3(\FIFO[103][23] ), .IN4(n6601), 
        .Q(n1258) );
  AO22X1 U2696 ( .IN1(n7096), .IN2(n6593), .IN3(\FIFO[102][0] ), .IN4(n6594), 
        .Q(n1267) );
  AO22X1 U2697 ( .IN1(n7068), .IN2(n6591), .IN3(\FIFO[102][2] ), .IN4(n6594), 
        .Q(n1269) );
  AO22X1 U2698 ( .IN1(n7057), .IN2(n6593), .IN3(\FIFO[102][3] ), .IN4(n6594), 
        .Q(n1270) );
  AO22X1 U2699 ( .IN1(n7046), .IN2(n6592), .IN3(\FIFO[102][4] ), .IN4(n6594), 
        .Q(n1271) );
  AO22X1 U2700 ( .IN1(n7035), .IN2(n6591), .IN3(\FIFO[102][5] ), .IN4(n6594), 
        .Q(n1272) );
  AO22X1 U2701 ( .IN1(n7024), .IN2(n6593), .IN3(\FIFO[102][6] ), .IN4(n6594), 
        .Q(n1273) );
  AO22X1 U2702 ( .IN1(n7013), .IN2(n6593), .IN3(\FIFO[102][7] ), .IN4(n6594), 
        .Q(n1274) );
  AO22X1 U2703 ( .IN1(n7002), .IN2(n6593), .IN3(\FIFO[102][8] ), .IN4(n6594), 
        .Q(n1275) );
  AO22X1 U2704 ( .IN1(n6991), .IN2(n6593), .IN3(\FIFO[102][9] ), .IN4(n6594), 
        .Q(n1276) );
  AO22X1 U2705 ( .IN1(n6980), .IN2(n6593), .IN3(\FIFO[102][10] ), .IN4(n6594), 
        .Q(n1277) );
  AO22X1 U2706 ( .IN1(n6969), .IN2(n6593), .IN3(\FIFO[102][11] ), .IN4(n6594), 
        .Q(n1278) );
  AO22X1 U2707 ( .IN1(n6958), .IN2(n6593), .IN3(\FIFO[102][12] ), .IN4(n6595), 
        .Q(n1279) );
  AO22X1 U2708 ( .IN1(n6947), .IN2(n6593), .IN3(\FIFO[102][13] ), .IN4(n6595), 
        .Q(n1280) );
  AO22X1 U2709 ( .IN1(n6936), .IN2(n6592), .IN3(\FIFO[102][14] ), .IN4(n6595), 
        .Q(n1281) );
  AO22X1 U2710 ( .IN1(n6925), .IN2(n6592), .IN3(\FIFO[102][15] ), .IN4(n6595), 
        .Q(n1282) );
  AO22X1 U2711 ( .IN1(n6914), .IN2(n6592), .IN3(\FIFO[102][16] ), .IN4(n6595), 
        .Q(n1283) );
  AO22X1 U2712 ( .IN1(n6903), .IN2(n6592), .IN3(\FIFO[102][17] ), .IN4(n6595), 
        .Q(n1284) );
  AO22X1 U2713 ( .IN1(n6892), .IN2(n6592), .IN3(\FIFO[102][18] ), .IN4(n6595), 
        .Q(n1285) );
  AO22X1 U2714 ( .IN1(n6881), .IN2(n6592), .IN3(\FIFO[102][19] ), .IN4(n6595), 
        .Q(n1286) );
  AO22X1 U2715 ( .IN1(n6870), .IN2(n6592), .IN3(\FIFO[102][20] ), .IN4(n6595), 
        .Q(n1287) );
  AO22X1 U2716 ( .IN1(n6859), .IN2(n6591), .IN3(\FIFO[102][21] ), .IN4(n6595), 
        .Q(n1288) );
  AO22X1 U2717 ( .IN1(n6848), .IN2(n6591), .IN3(\FIFO[102][22] ), .IN4(n6595), 
        .Q(n1289) );
  AO22X1 U2718 ( .IN1(n6837), .IN2(n6591), .IN3(\FIFO[102][23] ), .IN4(n6595), 
        .Q(n1290) );
  AO22X1 U2746 ( .IN1(n7096), .IN2(n6575), .IN3(\FIFO[99][0] ), .IN4(n6576), 
        .Q(n1363) );
  AO22X1 U2766 ( .IN1(n7079), .IN2(n6575), .IN3(\FIFO[99][1] ), .IN4(n6576), 
        .Q(n1364) );
  AO22X1 U2780 ( .IN1(n7068), .IN2(n6575), .IN3(\FIFO[99][2] ), .IN4(n6576), 
        .Q(n1365) );
  AO22X1 U2794 ( .IN1(n7057), .IN2(n6575), .IN3(\FIFO[99][3] ), .IN4(n6576), 
        .Q(n1366) );
  AO22X1 U2795 ( .IN1(n7046), .IN2(n6575), .IN3(\FIFO[99][4] ), .IN4(n6576), 
        .Q(n1367) );
  AO22X1 U2796 ( .IN1(n7035), .IN2(n6575), .IN3(\FIFO[99][5] ), .IN4(n6576), 
        .Q(n1368) );
  AO22X1 U2797 ( .IN1(n7024), .IN2(n6575), .IN3(\FIFO[99][6] ), .IN4(n6576), 
        .Q(n1369) );
  AO22X1 U2798 ( .IN1(n7013), .IN2(n6574), .IN3(\FIFO[99][7] ), .IN4(n6576), 
        .Q(n1370) );
  AO22X1 U2799 ( .IN1(n7002), .IN2(n6574), .IN3(\FIFO[99][8] ), .IN4(n6576), 
        .Q(n1371) );
  AO22X1 U2800 ( .IN1(n6991), .IN2(n6574), .IN3(\FIFO[99][9] ), .IN4(n6576), 
        .Q(n1372) );
  AO22X1 U2801 ( .IN1(n6980), .IN2(n6574), .IN3(\FIFO[99][10] ), .IN4(n6576), 
        .Q(n1373) );
  AO22X1 U2802 ( .IN1(n6969), .IN2(n6574), .IN3(\FIFO[99][11] ), .IN4(n6576), 
        .Q(n1374) );
  AO22X1 U2803 ( .IN1(n6958), .IN2(n6574), .IN3(\FIFO[99][12] ), .IN4(n6577), 
        .Q(n1375) );
  AO22X1 U2804 ( .IN1(n6947), .IN2(n6574), .IN3(\FIFO[99][13] ), .IN4(n6577), 
        .Q(n1376) );
  AO22X1 U2805 ( .IN1(n6936), .IN2(n6573), .IN3(\FIFO[99][14] ), .IN4(n6577), 
        .Q(n1377) );
  AO22X1 U2806 ( .IN1(n6925), .IN2(n6573), .IN3(\FIFO[99][15] ), .IN4(n6577), 
        .Q(n1378) );
  AO22X1 U2807 ( .IN1(n6914), .IN2(n6573), .IN3(\FIFO[99][16] ), .IN4(n6577), 
        .Q(n1379) );
  AO22X1 U2808 ( .IN1(n6903), .IN2(n6573), .IN3(\FIFO[99][17] ), .IN4(n6577), 
        .Q(n1380) );
  AO22X1 U2809 ( .IN1(n6892), .IN2(n6573), .IN3(\FIFO[99][18] ), .IN4(n6577), 
        .Q(n1381) );
  AO22X1 U2810 ( .IN1(n6881), .IN2(n6573), .IN3(\FIFO[99][19] ), .IN4(n6577), 
        .Q(n1382) );
  AO22X1 U2811 ( .IN1(n6870), .IN2(n6573), .IN3(\FIFO[99][20] ), .IN4(n6577), 
        .Q(n1383) );
  AO22X1 U2812 ( .IN1(n6859), .IN2(n6575), .IN3(\FIFO[99][21] ), .IN4(n6577), 
        .Q(n1384) );
  AO22X1 U2813 ( .IN1(n6848), .IN2(n6574), .IN3(\FIFO[99][22] ), .IN4(n6577), 
        .Q(n1385) );
  AO22X1 U2814 ( .IN1(n6837), .IN2(n6573), .IN3(\FIFO[99][23] ), .IN4(n6577), 
        .Q(n1386) );
  AO22X1 U2815 ( .IN1(n7096), .IN2(n6569), .IN3(\FIFO[98][0] ), .IN4(n6570), 
        .Q(n1395) );
  AO22X1 U2816 ( .IN1(n7079), .IN2(n6569), .IN3(\FIFO[98][1] ), .IN4(n6570), 
        .Q(n1396) );
  AO22X1 U2817 ( .IN1(n7068), .IN2(n6569), .IN3(\FIFO[98][2] ), .IN4(n6570), 
        .Q(n1397) );
  AO22X1 U2827 ( .IN1(n7057), .IN2(n6569), .IN3(\FIFO[98][3] ), .IN4(n6570), 
        .Q(n1398) );
  AO22X1 U2828 ( .IN1(n7046), .IN2(n6569), .IN3(\FIFO[98][4] ), .IN4(n6570), 
        .Q(n1399) );
  AO22X1 U2829 ( .IN1(n7035), .IN2(n6569), .IN3(\FIFO[98][5] ), .IN4(n6570), 
        .Q(n1400) );
  AO22X1 U2830 ( .IN1(n7024), .IN2(n6569), .IN3(\FIFO[98][6] ), .IN4(n6570), 
        .Q(n1401) );
  AO22X1 U2831 ( .IN1(n7013), .IN2(n6568), .IN3(\FIFO[98][7] ), .IN4(n6570), 
        .Q(n1402) );
  AO22X1 U2832 ( .IN1(n7002), .IN2(n6568), .IN3(\FIFO[98][8] ), .IN4(n6570), 
        .Q(n1403) );
  AO22X1 U2833 ( .IN1(n6991), .IN2(n6568), .IN3(\FIFO[98][9] ), .IN4(n6570), 
        .Q(n1404) );
  AO22X1 U2834 ( .IN1(n6980), .IN2(n6568), .IN3(\FIFO[98][10] ), .IN4(n6570), 
        .Q(n1405) );
  AO22X1 U2835 ( .IN1(n6969), .IN2(n6568), .IN3(\FIFO[98][11] ), .IN4(n6570), 
        .Q(n1406) );
  AO22X1 U2836 ( .IN1(n6958), .IN2(n6568), .IN3(\FIFO[98][12] ), .IN4(n6571), 
        .Q(n1407) );
  AO22X1 U2837 ( .IN1(n6936), .IN2(n6569), .IN3(\FIFO[98][14] ), .IN4(n6571), 
        .Q(n1409) );
  AO22X1 U2838 ( .IN1(n6925), .IN2(n6568), .IN3(\FIFO[98][15] ), .IN4(n6571), 
        .Q(n1410) );
  AO22X1 U2839 ( .IN1(n6914), .IN2(n6567), .IN3(\FIFO[98][16] ), .IN4(n6571), 
        .Q(n1411) );
  AO22X1 U2840 ( .IN1(n6903), .IN2(n6569), .IN3(\FIFO[98][17] ), .IN4(n6571), 
        .Q(n1412) );
  AO22X1 U2841 ( .IN1(n6892), .IN2(n6568), .IN3(\FIFO[98][18] ), .IN4(n6571), 
        .Q(n1413) );
  AO22X1 U2842 ( .IN1(n6881), .IN2(n6567), .IN3(\FIFO[98][19] ), .IN4(n6571), 
        .Q(n1414) );
  AO22X1 U2843 ( .IN1(n6870), .IN2(n6569), .IN3(\FIFO[98][20] ), .IN4(n6571), 
        .Q(n1415) );
  AO22X1 U2844 ( .IN1(n6859), .IN2(n6567), .IN3(\FIFO[98][21] ), .IN4(n6571), 
        .Q(n1416) );
  AO22X1 U2845 ( .IN1(n6848), .IN2(n6567), .IN3(\FIFO[98][22] ), .IN4(n6571), 
        .Q(n1417) );
  AO22X1 U2846 ( .IN1(n6837), .IN2(n6567), .IN3(\FIFO[98][23] ), .IN4(n6571), 
        .Q(n1418) );
  AO22X1 U2847 ( .IN1(n7095), .IN2(n6551), .IN3(\FIFO[95][0] ), .IN4(n6552), 
        .Q(n1491) );
  AO22X1 U2848 ( .IN1(n7078), .IN2(n6551), .IN3(\FIFO[95][1] ), .IN4(n6552), 
        .Q(n1492) );
  AO22X1 U2849 ( .IN1(n7067), .IN2(n6551), .IN3(\FIFO[95][2] ), .IN4(n6552), 
        .Q(n1493) );
  AO22X1 U2850 ( .IN1(n7056), .IN2(n6551), .IN3(\FIFO[95][3] ), .IN4(n6552), 
        .Q(n1494) );
  AO22X1 U2904 ( .IN1(n7045), .IN2(n6551), .IN3(\FIFO[95][4] ), .IN4(n6552), 
        .Q(n1495) );
  AO22X1 U2913 ( .IN1(n7034), .IN2(n6551), .IN3(\FIFO[95][5] ), .IN4(n6552), 
        .Q(n1496) );
  AO22X1 U2926 ( .IN1(n7023), .IN2(n6551), .IN3(\FIFO[95][6] ), .IN4(n6552), 
        .Q(n1497) );
  AO22X1 U2927 ( .IN1(n7012), .IN2(n6550), .IN3(\FIFO[95][7] ), .IN4(n6552), 
        .Q(n1498) );
  AO22X1 U2928 ( .IN1(n7001), .IN2(n6550), .IN3(\FIFO[95][8] ), .IN4(n6552), 
        .Q(n1499) );
  AO22X1 U2929 ( .IN1(n6990), .IN2(n6550), .IN3(\FIFO[95][9] ), .IN4(n6552), 
        .Q(n1500) );
  AO22X1 U2930 ( .IN1(n6979), .IN2(n6550), .IN3(\FIFO[95][10] ), .IN4(n6552), 
        .Q(n1501) );
  AO22X1 U2931 ( .IN1(n6968), .IN2(n6550), .IN3(\FIFO[95][11] ), .IN4(n6552), 
        .Q(n1502) );
  AO22X1 U2932 ( .IN1(n6957), .IN2(n6550), .IN3(\FIFO[95][12] ), .IN4(n6553), 
        .Q(n1503) );
  AO22X1 U2933 ( .IN1(n6946), .IN2(n6550), .IN3(\FIFO[95][13] ), .IN4(n6553), 
        .Q(n1504) );
  AO22X1 U2934 ( .IN1(n6935), .IN2(n6549), .IN3(\FIFO[95][14] ), .IN4(n6553), 
        .Q(n1505) );
  AO22X1 U2935 ( .IN1(n6924), .IN2(n6549), .IN3(\FIFO[95][15] ), .IN4(n6553), 
        .Q(n1506) );
  AO22X1 U2936 ( .IN1(n6913), .IN2(n6549), .IN3(\FIFO[95][16] ), .IN4(n6553), 
        .Q(n1507) );
  AO22X1 U2937 ( .IN1(n6902), .IN2(n6549), .IN3(\FIFO[95][17] ), .IN4(n6553), 
        .Q(n1508) );
  AO22X1 U2938 ( .IN1(n6891), .IN2(n6549), .IN3(\FIFO[95][18] ), .IN4(n6553), 
        .Q(n1509) );
  AO22X1 U2939 ( .IN1(n6880), .IN2(n6549), .IN3(\FIFO[95][19] ), .IN4(n6553), 
        .Q(n1510) );
  AO22X1 U2940 ( .IN1(n6869), .IN2(n6549), .IN3(\FIFO[95][20] ), .IN4(n6553), 
        .Q(n1511) );
  AO22X1 U2941 ( .IN1(n6858), .IN2(n6551), .IN3(\FIFO[95][21] ), .IN4(n6553), 
        .Q(n1512) );
  AO22X1 U2942 ( .IN1(n6847), .IN2(n6550), .IN3(\FIFO[95][22] ), .IN4(n6553), 
        .Q(n1513) );
  AO22X1 U2943 ( .IN1(n6836), .IN2(n6549), .IN3(\FIFO[95][23] ), .IN4(n6553), 
        .Q(n1514) );
  AO22X1 U2944 ( .IN1(n7095), .IN2(n6545), .IN3(\FIFO[94][0] ), .IN4(n6546), 
        .Q(n1523) );
  AO22X1 U2945 ( .IN1(n7067), .IN2(n6545), .IN3(\FIFO[94][2] ), .IN4(n6546), 
        .Q(n1525) );
  AO22X1 U2946 ( .IN1(n7056), .IN2(n6545), .IN3(\FIFO[94][3] ), .IN4(n6546), 
        .Q(n1526) );
  AO22X1 U2947 ( .IN1(n7045), .IN2(n6545), .IN3(\FIFO[94][4] ), .IN4(n6546), 
        .Q(n1527) );
  AO22X1 U2948 ( .IN1(n7034), .IN2(n6545), .IN3(\FIFO[94][5] ), .IN4(n6546), 
        .Q(n1528) );
  AO22X1 U2949 ( .IN1(n7023), .IN2(n6545), .IN3(\FIFO[94][6] ), .IN4(n6546), 
        .Q(n1529) );
  AO22X1 U2950 ( .IN1(n7012), .IN2(n6544), .IN3(\FIFO[94][7] ), .IN4(n6546), 
        .Q(n1530) );
  AO22X1 U2960 ( .IN1(n7001), .IN2(n6544), .IN3(\FIFO[94][8] ), .IN4(n6546), 
        .Q(n1531) );
  AO22X1 U2961 ( .IN1(n6990), .IN2(n6544), .IN3(\FIFO[94][9] ), .IN4(n6546), 
        .Q(n1532) );
  AO22X1 U2962 ( .IN1(n6979), .IN2(n6544), .IN3(\FIFO[94][10] ), .IN4(n6546), 
        .Q(n1533) );
  AO22X1 U2963 ( .IN1(n6968), .IN2(n6544), .IN3(\FIFO[94][11] ), .IN4(n6546), 
        .Q(n1534) );
  AO22X1 U2964 ( .IN1(n6957), .IN2(n6544), .IN3(\FIFO[94][12] ), .IN4(n6547), 
        .Q(n1535) );
  AO22X1 U2965 ( .IN1(n6946), .IN2(n6544), .IN3(\FIFO[94][13] ), .IN4(n6547), 
        .Q(n1536) );
  AO22X1 U2966 ( .IN1(n6935), .IN2(n6545), .IN3(\FIFO[94][14] ), .IN4(n6547), 
        .Q(n1537) );
  AO22X1 U2967 ( .IN1(n6913), .IN2(n6543), .IN3(\FIFO[94][16] ), .IN4(n6547), 
        .Q(n1539) );
  AO22X1 U2968 ( .IN1(n6902), .IN2(n6545), .IN3(\FIFO[94][17] ), .IN4(n6547), 
        .Q(n1540) );
  AO22X1 U2969 ( .IN1(n6891), .IN2(n6544), .IN3(\FIFO[94][18] ), .IN4(n6547), 
        .Q(n1541) );
  AO22X1 U2970 ( .IN1(n6880), .IN2(n6543), .IN3(\FIFO[94][19] ), .IN4(n6547), 
        .Q(n1542) );
  AO22X1 U2971 ( .IN1(n6869), .IN2(n6545), .IN3(\FIFO[94][20] ), .IN4(n6547), 
        .Q(n1543) );
  AO22X1 U2972 ( .IN1(n6858), .IN2(n6543), .IN3(\FIFO[94][21] ), .IN4(n6547), 
        .Q(n1544) );
  AO22X1 U2973 ( .IN1(n6847), .IN2(n6543), .IN3(\FIFO[94][22] ), .IN4(n6547), 
        .Q(n1545) );
  AO22X1 U2974 ( .IN1(n6836), .IN2(n6543), .IN3(\FIFO[94][23] ), .IN4(n6547), 
        .Q(n1546) );
  AO22X1 U2975 ( .IN1(n7095), .IN2(n6527), .IN3(\FIFO[91][0] ), .IN4(n6528), 
        .Q(n1619) );
  AO22X1 U2976 ( .IN1(n7078), .IN2(n6527), .IN3(\FIFO[91][1] ), .IN4(n6528), 
        .Q(n1620) );
  AO22X1 U2977 ( .IN1(n7067), .IN2(n6527), .IN3(\FIFO[91][2] ), .IN4(n6528), 
        .Q(n1621) );
  AO22X1 U2978 ( .IN1(n7056), .IN2(n6527), .IN3(\FIFO[91][3] ), .IN4(n6528), 
        .Q(n1622) );
  AO22X1 U2979 ( .IN1(n7045), .IN2(n6527), .IN3(\FIFO[91][4] ), .IN4(n6528), 
        .Q(n1623) );
  AO22X1 U2980 ( .IN1(n7034), .IN2(n6527), .IN3(\FIFO[91][5] ), .IN4(n6528), 
        .Q(n1624) );
  AO22X1 U2981 ( .IN1(n7023), .IN2(n6527), .IN3(\FIFO[91][6] ), .IN4(n6528), 
        .Q(n1625) );
  AO22X1 U2982 ( .IN1(n7012), .IN2(n6526), .IN3(\FIFO[91][7] ), .IN4(n6528), 
        .Q(n1626) );
  AO22X1 U2983 ( .IN1(n7001), .IN2(n6526), .IN3(\FIFO[91][8] ), .IN4(n6528), 
        .Q(n1627) );
  AO22X1 U3026 ( .IN1(n6990), .IN2(n6526), .IN3(\FIFO[91][9] ), .IN4(n6528), 
        .Q(n1628) );
  AO22X1 U3047 ( .IN1(n6979), .IN2(n6526), .IN3(\FIFO[91][10] ), .IN4(n6528), 
        .Q(n1629) );
  AO22X1 U3059 ( .IN1(n6968), .IN2(n6526), .IN3(\FIFO[91][11] ), .IN4(n6528), 
        .Q(n1630) );
  AO22X1 U3060 ( .IN1(n6957), .IN2(n6526), .IN3(\FIFO[91][12] ), .IN4(n6529), 
        .Q(n1631) );
  AO22X1 U3061 ( .IN1(n6946), .IN2(n6526), .IN3(\FIFO[91][13] ), .IN4(n6529), 
        .Q(n1632) );
  AO22X1 U3062 ( .IN1(n6935), .IN2(n6525), .IN3(\FIFO[91][14] ), .IN4(n6529), 
        .Q(n1633) );
  AO22X1 U3063 ( .IN1(n6924), .IN2(n6525), .IN3(\FIFO[91][15] ), .IN4(n6529), 
        .Q(n1634) );
  AO22X1 U3064 ( .IN1(n6913), .IN2(n6525), .IN3(\FIFO[91][16] ), .IN4(n6529), 
        .Q(n1635) );
  AO22X1 U3065 ( .IN1(n6902), .IN2(n6525), .IN3(\FIFO[91][17] ), .IN4(n6529), 
        .Q(n1636) );
  AO22X1 U3066 ( .IN1(n6891), .IN2(n6525), .IN3(\FIFO[91][18] ), .IN4(n6529), 
        .Q(n1637) );
  AO22X1 U3067 ( .IN1(n6880), .IN2(n6525), .IN3(\FIFO[91][19] ), .IN4(n6529), 
        .Q(n1638) );
  AO22X1 U3068 ( .IN1(n6869), .IN2(n6525), .IN3(\FIFO[91][20] ), .IN4(n6529), 
        .Q(n1639) );
  AO22X1 U3069 ( .IN1(n6858), .IN2(n6527), .IN3(\FIFO[91][21] ), .IN4(n6529), 
        .Q(n1640) );
  AO22X1 U3070 ( .IN1(n6847), .IN2(n6526), .IN3(\FIFO[91][22] ), .IN4(n6529), 
        .Q(n1641) );
  AO22X1 U3071 ( .IN1(n6836), .IN2(n6525), .IN3(\FIFO[91][23] ), .IN4(n6529), 
        .Q(n1642) );
  AO22X1 U3072 ( .IN1(n7095), .IN2(n6521), .IN3(\FIFO[90][0] ), .IN4(n6522), 
        .Q(n1651) );
  AO22X1 U3073 ( .IN1(n7078), .IN2(n6521), .IN3(\FIFO[90][1] ), .IN4(n6522), 
        .Q(n1652) );
  AO22X1 U3074 ( .IN1(n7067), .IN2(n6521), .IN3(\FIFO[90][2] ), .IN4(n6522), 
        .Q(n1653) );
  AO22X1 U3075 ( .IN1(n7056), .IN2(n6521), .IN3(\FIFO[90][3] ), .IN4(n6522), 
        .Q(n1654) );
  AO22X1 U3076 ( .IN1(n7045), .IN2(n6521), .IN3(\FIFO[90][4] ), .IN4(n6522), 
        .Q(n1655) );
  AO22X1 U3077 ( .IN1(n7034), .IN2(n6521), .IN3(\FIFO[90][5] ), .IN4(n6522), 
        .Q(n1656) );
  AO22X1 U3078 ( .IN1(n7023), .IN2(n6521), .IN3(\FIFO[90][6] ), .IN4(n6522), 
        .Q(n1657) );
  AO22X1 U3079 ( .IN1(n7012), .IN2(n6520), .IN3(\FIFO[90][7] ), .IN4(n6522), 
        .Q(n1658) );
  AO22X1 U3080 ( .IN1(n7001), .IN2(n6520), .IN3(\FIFO[90][8] ), .IN4(n6522), 
        .Q(n1659) );
  AO22X1 U3081 ( .IN1(n6990), .IN2(n6520), .IN3(\FIFO[90][9] ), .IN4(n6522), 
        .Q(n1660) );
  AO22X1 U3082 ( .IN1(n6979), .IN2(n6520), .IN3(\FIFO[90][10] ), .IN4(n6522), 
        .Q(n1661) );
  AO22X1 U3092 ( .IN1(n6968), .IN2(n6520), .IN3(\FIFO[90][11] ), .IN4(n6522), 
        .Q(n1662) );
  AO22X1 U3093 ( .IN1(n6957), .IN2(n6520), .IN3(\FIFO[90][12] ), .IN4(n6523), 
        .Q(n1663) );
  AO22X1 U3094 ( .IN1(n6946), .IN2(n6520), .IN3(\FIFO[90][13] ), .IN4(n6523), 
        .Q(n1664) );
  AO22X1 U3095 ( .IN1(n6935), .IN2(n6519), .IN3(\FIFO[90][14] ), .IN4(n6523), 
        .Q(n1665) );
  AO22X1 U3096 ( .IN1(n6924), .IN2(n6519), .IN3(\FIFO[90][15] ), .IN4(n6523), 
        .Q(n1666) );
  AO22X1 U3097 ( .IN1(n6913), .IN2(n6519), .IN3(\FIFO[90][16] ), .IN4(n6523), 
        .Q(n1667) );
  AO22X1 U3098 ( .IN1(n6902), .IN2(n6519), .IN3(\FIFO[90][17] ), .IN4(n6523), 
        .Q(n1668) );
  AO22X1 U3099 ( .IN1(n6891), .IN2(n6519), .IN3(\FIFO[90][18] ), .IN4(n6523), 
        .Q(n1669) );
  AO22X1 U3100 ( .IN1(n6880), .IN2(n6519), .IN3(\FIFO[90][19] ), .IN4(n6523), 
        .Q(n1670) );
  AO22X1 U3101 ( .IN1(n6869), .IN2(n6519), .IN3(\FIFO[90][20] ), .IN4(n6523), 
        .Q(n1671) );
  AO22X1 U3102 ( .IN1(n6858), .IN2(n6521), .IN3(\FIFO[90][21] ), .IN4(n6523), 
        .Q(n1672) );
  AO22X1 U3103 ( .IN1(n6847), .IN2(n6520), .IN3(\FIFO[90][22] ), .IN4(n6523), 
        .Q(n1673) );
  AO22X1 U3104 ( .IN1(n6836), .IN2(n6519), .IN3(\FIFO[90][23] ), .IN4(n6523), 
        .Q(n1674) );
  AO22X1 U3105 ( .IN1(n7095), .IN2(n6503), .IN3(\FIFO[87][0] ), .IN4(n6504), 
        .Q(n1747) );
  AO22X1 U3106 ( .IN1(n7078), .IN2(n6503), .IN3(\FIFO[87][1] ), .IN4(n6504), 
        .Q(n1748) );
  AO22X1 U3107 ( .IN1(n7067), .IN2(n6503), .IN3(\FIFO[87][2] ), .IN4(n6504), 
        .Q(n1749) );
  AO22X1 U3108 ( .IN1(n7056), .IN2(n6503), .IN3(\FIFO[87][3] ), .IN4(n6504), 
        .Q(n1750) );
  AO22X1 U3109 ( .IN1(n7045), .IN2(n6503), .IN3(\FIFO[87][4] ), .IN4(n6504), 
        .Q(n1751) );
  AO22X1 U3110 ( .IN1(n7034), .IN2(n6503), .IN3(\FIFO[87][5] ), .IN4(n6504), 
        .Q(n1752) );
  AO22X1 U3111 ( .IN1(n7023), .IN2(n6503), .IN3(\FIFO[87][6] ), .IN4(n6504), 
        .Q(n1753) );
  AO22X1 U3112 ( .IN1(n7012), .IN2(n6502), .IN3(\FIFO[87][7] ), .IN4(n6504), 
        .Q(n1754) );
  AO22X1 U3113 ( .IN1(n7001), .IN2(n6502), .IN3(\FIFO[87][8] ), .IN4(n6504), 
        .Q(n1755) );
  AO22X1 U3114 ( .IN1(n6990), .IN2(n6502), .IN3(\FIFO[87][9] ), .IN4(n6504), 
        .Q(n1756) );
  AO22X1 U3115 ( .IN1(n6979), .IN2(n6502), .IN3(\FIFO[87][10] ), .IN4(n6504), 
        .Q(n1757) );
  AO22X1 U3133 ( .IN1(n6968), .IN2(n6502), .IN3(\FIFO[87][11] ), .IN4(n6504), 
        .Q(n1758) );
  AO22X1 U3167 ( .IN1(n6957), .IN2(n6502), .IN3(\FIFO[87][12] ), .IN4(n6505), 
        .Q(n1759) );
  AO22X1 U3191 ( .IN1(n6946), .IN2(n6502), .IN3(\FIFO[87][13] ), .IN4(n6505), 
        .Q(n1760) );
  AO22X1 U3192 ( .IN1(n6935), .IN2(n6501), .IN3(\FIFO[87][14] ), .IN4(n6505), 
        .Q(n1761) );
  AO22X1 U3193 ( .IN1(n6924), .IN2(n6501), .IN3(\FIFO[87][15] ), .IN4(n6505), 
        .Q(n1762) );
  AO22X1 U3194 ( .IN1(n6913), .IN2(n6501), .IN3(\FIFO[87][16] ), .IN4(n6505), 
        .Q(n1763) );
  AO22X1 U3195 ( .IN1(n6902), .IN2(n6501), .IN3(\FIFO[87][17] ), .IN4(n6505), 
        .Q(n1764) );
  AO22X1 U3196 ( .IN1(n6891), .IN2(n6501), .IN3(\FIFO[87][18] ), .IN4(n6505), 
        .Q(n1765) );
  AO22X1 U3197 ( .IN1(n6880), .IN2(n6501), .IN3(\FIFO[87][19] ), .IN4(n6505), 
        .Q(n1766) );
  AO22X1 U3198 ( .IN1(n6869), .IN2(n6501), .IN3(\FIFO[87][20] ), .IN4(n6505), 
        .Q(n1767) );
  AO22X1 U3199 ( .IN1(n6858), .IN2(n6503), .IN3(\FIFO[87][21] ), .IN4(n6505), 
        .Q(n1768) );
  AO22X1 U3200 ( .IN1(n6847), .IN2(n6502), .IN3(\FIFO[87][22] ), .IN4(n6505), 
        .Q(n1769) );
  AO22X1 U3201 ( .IN1(n6836), .IN2(n6501), .IN3(\FIFO[87][23] ), .IN4(n6505), 
        .Q(n1770) );
  AO22X1 U3202 ( .IN1(n7095), .IN2(n6497), .IN3(\FIFO[86][0] ), .IN4(n6498), 
        .Q(n1779) );
  AO22X1 U3203 ( .IN1(n7078), .IN2(n6497), .IN3(\FIFO[86][1] ), .IN4(n6498), 
        .Q(n1780) );
  AO22X1 U3204 ( .IN1(n7067), .IN2(n6497), .IN3(\FIFO[86][2] ), .IN4(n6498), 
        .Q(n1781) );
  AO22X1 U3205 ( .IN1(n7056), .IN2(n6497), .IN3(\FIFO[86][3] ), .IN4(n6498), 
        .Q(n1782) );
  AO22X1 U3206 ( .IN1(n7045), .IN2(n6497), .IN3(\FIFO[86][4] ), .IN4(n6498), 
        .Q(n1783) );
  AO22X1 U3207 ( .IN1(n7034), .IN2(n6497), .IN3(\FIFO[86][5] ), .IN4(n6498), 
        .Q(n1784) );
  AO22X1 U3208 ( .IN1(n7023), .IN2(n6497), .IN3(\FIFO[86][6] ), .IN4(n6498), 
        .Q(n1785) );
  AO22X1 U3209 ( .IN1(n7012), .IN2(n6496), .IN3(\FIFO[86][7] ), .IN4(n6498), 
        .Q(n1786) );
  AO22X1 U3210 ( .IN1(n7001), .IN2(n6496), .IN3(\FIFO[86][8] ), .IN4(n6498), 
        .Q(n1787) );
  AO22X1 U3211 ( .IN1(n6990), .IN2(n6496), .IN3(\FIFO[86][9] ), .IN4(n6498), 
        .Q(n1788) );
  AO22X1 U3212 ( .IN1(n6979), .IN2(n6496), .IN3(\FIFO[86][10] ), .IN4(n6498), 
        .Q(n1789) );
  AO22X1 U3213 ( .IN1(n6968), .IN2(n6496), .IN3(\FIFO[86][11] ), .IN4(n6498), 
        .Q(n1790) );
  AO22X1 U3214 ( .IN1(n6957), .IN2(n6496), .IN3(\FIFO[86][12] ), .IN4(n6499), 
        .Q(n1791) );
  AO22X1 U3224 ( .IN1(n6946), .IN2(n6496), .IN3(\FIFO[86][13] ), .IN4(n6499), 
        .Q(n1792) );
  AO22X1 U3225 ( .IN1(n6935), .IN2(n6495), .IN3(\FIFO[86][14] ), .IN4(n6499), 
        .Q(n1793) );
  AO22X1 U3226 ( .IN1(n6924), .IN2(n6495), .IN3(\FIFO[86][15] ), .IN4(n6499), 
        .Q(n1794) );
  AO22X1 U3227 ( .IN1(n6913), .IN2(n6495), .IN3(\FIFO[86][16] ), .IN4(n6499), 
        .Q(n1795) );
  AO22X1 U3228 ( .IN1(n6902), .IN2(n6495), .IN3(\FIFO[86][17] ), .IN4(n6499), 
        .Q(n1796) );
  AO22X1 U3229 ( .IN1(n6891), .IN2(n6495), .IN3(\FIFO[86][18] ), .IN4(n6499), 
        .Q(n1797) );
  AO22X1 U3230 ( .IN1(n6880), .IN2(n6495), .IN3(\FIFO[86][19] ), .IN4(n6499), 
        .Q(n1798) );
  AO22X1 U3231 ( .IN1(n6869), .IN2(n6495), .IN3(\FIFO[86][20] ), .IN4(n6499), 
        .Q(n1799) );
  AO22X1 U3232 ( .IN1(n6858), .IN2(n6497), .IN3(\FIFO[86][21] ), .IN4(n6499), 
        .Q(n1800) );
  AO22X1 U3233 ( .IN1(n6847), .IN2(n6496), .IN3(\FIFO[86][22] ), .IN4(n6499), 
        .Q(n1801) );
  AO22X1 U3234 ( .IN1(n6836), .IN2(n6495), .IN3(\FIFO[86][23] ), .IN4(n6499), 
        .Q(n1802) );
  AO22X1 U3235 ( .IN1(n7094), .IN2(n6479), .IN3(\FIFO[83][0] ), .IN4(n6480), 
        .Q(n1875) );
  AO22X1 U3236 ( .IN1(n7077), .IN2(n6478), .IN3(\FIFO[83][1] ), .IN4(n6480), 
        .Q(n1876) );
  AO22X1 U3237 ( .IN1(n7066), .IN2(n6477), .IN3(\FIFO[83][2] ), .IN4(n6480), 
        .Q(n1877) );
  AO22X1 U3238 ( .IN1(n7055), .IN2(n6479), .IN3(\FIFO[83][3] ), .IN4(n6480), 
        .Q(n1878) );
  AO22X1 U3239 ( .IN1(n7044), .IN2(n6478), .IN3(\FIFO[83][4] ), .IN4(n6480), 
        .Q(n1879) );
  AO22X1 U3240 ( .IN1(n7033), .IN2(n6477), .IN3(\FIFO[83][5] ), .IN4(n6480), 
        .Q(n1880) );
  AO22X1 U3241 ( .IN1(n7011), .IN2(n6479), .IN3(\FIFO[83][7] ), .IN4(n6480), 
        .Q(n1882) );
  AO22X1 U3242 ( .IN1(n7000), .IN2(n6479), .IN3(\FIFO[83][8] ), .IN4(n6480), 
        .Q(n1883) );
  AO22X1 U3243 ( .IN1(n6989), .IN2(n6479), .IN3(\FIFO[83][9] ), .IN4(n6480), 
        .Q(n1884) );
  AO22X1 U3244 ( .IN1(n6978), .IN2(n6479), .IN3(\FIFO[83][10] ), .IN4(n6480), 
        .Q(n1885) );
  AO22X1 U3245 ( .IN1(n6967), .IN2(n6479), .IN3(\FIFO[83][11] ), .IN4(n6480), 
        .Q(n1886) );
  AO22X1 U3246 ( .IN1(n6956), .IN2(n6479), .IN3(\FIFO[83][12] ), .IN4(n6481), 
        .Q(n1887) );
  AO22X1 U3247 ( .IN1(n6945), .IN2(n6479), .IN3(\FIFO[83][13] ), .IN4(n6481), 
        .Q(n1888) );
  AO22X1 U3248 ( .IN1(n6934), .IN2(n6478), .IN3(\FIFO[83][14] ), .IN4(n6481), 
        .Q(n1889) );
  AO22X1 U3267 ( .IN1(n6923), .IN2(n6478), .IN3(\FIFO[83][15] ), .IN4(n6481), 
        .Q(n1890) );
  AO22X1 U3302 ( .IN1(n6912), .IN2(n6478), .IN3(\FIFO[83][16] ), .IN4(n6481), 
        .Q(n1891) );
  AO22X1 U3323 ( .IN1(n6901), .IN2(n6478), .IN3(\FIFO[83][17] ), .IN4(n6481), 
        .Q(n1892) );
  AO22X1 U3324 ( .IN1(n6890), .IN2(n6478), .IN3(\FIFO[83][18] ), .IN4(n6481), 
        .Q(n1893) );
  AO22X1 U3325 ( .IN1(n6879), .IN2(n6478), .IN3(\FIFO[83][19] ), .IN4(n6481), 
        .Q(n1894) );
  AO22X1 U3326 ( .IN1(n6857), .IN2(n6477), .IN3(\FIFO[83][21] ), .IN4(n6481), 
        .Q(n1896) );
  AO22X1 U3327 ( .IN1(n6846), .IN2(n6477), .IN3(\FIFO[83][22] ), .IN4(n6481), 
        .Q(n1897) );
  AO22X1 U3328 ( .IN1(n6835), .IN2(n6477), .IN3(\FIFO[83][23] ), .IN4(n6481), 
        .Q(n1898) );
  AO22X1 U3329 ( .IN1(n7094), .IN2(n6473), .IN3(\FIFO[82][0] ), .IN4(n6474), 
        .Q(n1907) );
  AO22X1 U3330 ( .IN1(n7077), .IN2(n6473), .IN3(\FIFO[82][1] ), .IN4(n6474), 
        .Q(n1908) );
  AO22X1 U3331 ( .IN1(n7066), .IN2(n6473), .IN3(\FIFO[82][2] ), .IN4(n6474), 
        .Q(n1909) );
  AO22X1 U3332 ( .IN1(n7055), .IN2(n6473), .IN3(\FIFO[82][3] ), .IN4(n6474), 
        .Q(n1910) );
  AO22X1 U3333 ( .IN1(n7044), .IN2(n6473), .IN3(\FIFO[82][4] ), .IN4(n6474), 
        .Q(n1911) );
  AO22X1 U3334 ( .IN1(n7033), .IN2(n6473), .IN3(\FIFO[82][5] ), .IN4(n6474), 
        .Q(n1912) );
  AO22X1 U3335 ( .IN1(n7022), .IN2(n6473), .IN3(\FIFO[82][6] ), .IN4(n6474), 
        .Q(n1913) );
  AO22X1 U3336 ( .IN1(n7011), .IN2(n6472), .IN3(\FIFO[82][7] ), .IN4(n6474), 
        .Q(n1914) );
  AO22X1 U3337 ( .IN1(n7000), .IN2(n6472), .IN3(\FIFO[82][8] ), .IN4(n6474), 
        .Q(n1915) );
  AO22X1 U3338 ( .IN1(n6989), .IN2(n6472), .IN3(\FIFO[82][9] ), .IN4(n6474), 
        .Q(n1916) );
  AO22X1 U3339 ( .IN1(n6978), .IN2(n6472), .IN3(\FIFO[82][10] ), .IN4(n6474), 
        .Q(n1917) );
  AO22X1 U3340 ( .IN1(n6967), .IN2(n6472), .IN3(\FIFO[82][11] ), .IN4(n6474), 
        .Q(n1918) );
  AO22X1 U3341 ( .IN1(n6956), .IN2(n6472), .IN3(\FIFO[82][12] ), .IN4(n6475), 
        .Q(n1919) );
  AO22X1 U3342 ( .IN1(n6945), .IN2(n6472), .IN3(\FIFO[82][13] ), .IN4(n6475), 
        .Q(n1920) );
  AO22X1 U3343 ( .IN1(n6934), .IN2(n6471), .IN3(\FIFO[82][14] ), .IN4(n6475), 
        .Q(n1921) );
  AO22X1 U3344 ( .IN1(n6923), .IN2(n6471), .IN3(\FIFO[82][15] ), .IN4(n6475), 
        .Q(n1922) );
  AO22X1 U3345 ( .IN1(n6912), .IN2(n6471), .IN3(\FIFO[82][16] ), .IN4(n6475), 
        .Q(n1923) );
  AO22X1 U3346 ( .IN1(n6901), .IN2(n6471), .IN3(\FIFO[82][17] ), .IN4(n6475), 
        .Q(n1924) );
  AO22X1 U3356 ( .IN1(n6890), .IN2(n6471), .IN3(\FIFO[82][18] ), .IN4(n6475), 
        .Q(n1925) );
  AO22X1 U3357 ( .IN1(n6879), .IN2(n6471), .IN3(\FIFO[82][19] ), .IN4(n6475), 
        .Q(n1926) );
  AO22X1 U3358 ( .IN1(n6868), .IN2(n6471), .IN3(\FIFO[82][20] ), .IN4(n6475), 
        .Q(n1927) );
  AO22X1 U3359 ( .IN1(n6857), .IN2(n6473), .IN3(\FIFO[82][21] ), .IN4(n6475), 
        .Q(n1928) );
  AO22X1 U3360 ( .IN1(n6846), .IN2(n6472), .IN3(\FIFO[82][22] ), .IN4(n6475), 
        .Q(n1929) );
  AO22X1 U3361 ( .IN1(n6835), .IN2(n6471), .IN3(\FIFO[82][23] ), .IN4(n6475), 
        .Q(n1930) );
  AO22X1 U3362 ( .IN1(n7094), .IN2(n6455), .IN3(\FIFO[79][0] ), .IN4(n6456), 
        .Q(n2003) );
  AO22X1 U3363 ( .IN1(n7077), .IN2(n6455), .IN3(\FIFO[79][1] ), .IN4(n6456), 
        .Q(n2004) );
  AO22X1 U3364 ( .IN1(n7066), .IN2(n6455), .IN3(\FIFO[79][2] ), .IN4(n6456), 
        .Q(n2005) );
  AO22X1 U3365 ( .IN1(n7055), .IN2(n6455), .IN3(\FIFO[79][3] ), .IN4(n6456), 
        .Q(n2006) );
  AO22X1 U3366 ( .IN1(n7044), .IN2(n6455), .IN3(\FIFO[79][4] ), .IN4(n6456), 
        .Q(n2007) );
  AO22X1 U3367 ( .IN1(n7033), .IN2(n6455), .IN3(\FIFO[79][5] ), .IN4(n6456), 
        .Q(n2008) );
  AO22X1 U3368 ( .IN1(n7022), .IN2(n6455), .IN3(\FIFO[79][6] ), .IN4(n6456), 
        .Q(n2009) );
  AO22X1 U3369 ( .IN1(n7011), .IN2(n6454), .IN3(\FIFO[79][7] ), .IN4(n6456), 
        .Q(n2010) );
  AO22X1 U3370 ( .IN1(n7000), .IN2(n6454), .IN3(\FIFO[79][8] ), .IN4(n6456), 
        .Q(n2011) );
  AO22X1 U3371 ( .IN1(n6989), .IN2(n6454), .IN3(\FIFO[79][9] ), .IN4(n6456), 
        .Q(n2012) );
  AO22X1 U3372 ( .IN1(n6978), .IN2(n6454), .IN3(\FIFO[79][10] ), .IN4(n6456), 
        .Q(n2013) );
  AO22X1 U3373 ( .IN1(n6967), .IN2(n6454), .IN3(\FIFO[79][11] ), .IN4(n6456), 
        .Q(n2014) );
  AO22X1 U3374 ( .IN1(n6956), .IN2(n6454), .IN3(\FIFO[79][12] ), .IN4(n6457), 
        .Q(n2015) );
  AO22X1 U3375 ( .IN1(n6945), .IN2(n6454), .IN3(\FIFO[79][13] ), .IN4(n6457), 
        .Q(n2016) );
  AO22X1 U3376 ( .IN1(n6934), .IN2(n6453), .IN3(\FIFO[79][14] ), .IN4(n6457), 
        .Q(n2017) );
  AO22X1 U3377 ( .IN1(n6923), .IN2(n6453), .IN3(\FIFO[79][15] ), .IN4(n6457), 
        .Q(n2018) );
  AO22X1 U3378 ( .IN1(n6912), .IN2(n6453), .IN3(\FIFO[79][16] ), .IN4(n6457), 
        .Q(n2019) );
  AO22X1 U3379 ( .IN1(n6901), .IN2(n6453), .IN3(\FIFO[79][17] ), .IN4(n6457), 
        .Q(n2020) );
  AO22X1 U3381 ( .IN1(n6890), .IN2(n6453), .IN3(\FIFO[79][18] ), .IN4(n6457), 
        .Q(n2021) );
  AO22X1 U3407 ( .IN1(n6879), .IN2(n6453), .IN3(\FIFO[79][19] ), .IN4(n6457), 
        .Q(n2022) );
  AO22X1 U3415 ( .IN1(n6868), .IN2(n6453), .IN3(\FIFO[79][20] ), .IN4(n6457), 
        .Q(n2023) );
  AO22X1 U3437 ( .IN1(n6857), .IN2(n6455), .IN3(\FIFO[79][21] ), .IN4(n6457), 
        .Q(n2024) );
  AO22X1 U3456 ( .IN1(n6846), .IN2(n6454), .IN3(\FIFO[79][22] ), .IN4(n6457), 
        .Q(n2025) );
  AO22X1 U3457 ( .IN1(n6835), .IN2(n6453), .IN3(\FIFO[79][23] ), .IN4(n6457), 
        .Q(n2026) );
  AO22X1 U3458 ( .IN1(n7094), .IN2(n6449), .IN3(\FIFO[78][0] ), .IN4(n6450), 
        .Q(n2035) );
  AO22X1 U3459 ( .IN1(n7077), .IN2(n6449), .IN3(\FIFO[78][1] ), .IN4(n6450), 
        .Q(n2036) );
  AO22X1 U3460 ( .IN1(n7066), .IN2(n6449), .IN3(\FIFO[78][2] ), .IN4(n6450), 
        .Q(n2037) );
  AO22X1 U3461 ( .IN1(n7055), .IN2(n6449), .IN3(\FIFO[78][3] ), .IN4(n6450), 
        .Q(n2038) );
  AO22X1 U3462 ( .IN1(n7044), .IN2(n6449), .IN3(\FIFO[78][4] ), .IN4(n6450), 
        .Q(n2039) );
  AO22X1 U3463 ( .IN1(n7033), .IN2(n6449), .IN3(\FIFO[78][5] ), .IN4(n6450), 
        .Q(n2040) );
  AO22X1 U3464 ( .IN1(n7022), .IN2(n6449), .IN3(\FIFO[78][6] ), .IN4(n6450), 
        .Q(n2041) );
  AO22X1 U3465 ( .IN1(n7011), .IN2(n6448), .IN3(\FIFO[78][7] ), .IN4(n6450), 
        .Q(n2042) );
  AO22X1 U3466 ( .IN1(n7000), .IN2(n6448), .IN3(\FIFO[78][8] ), .IN4(n6450), 
        .Q(n2043) );
  AO22X1 U3467 ( .IN1(n6989), .IN2(n6448), .IN3(\FIFO[78][9] ), .IN4(n6450), 
        .Q(n2044) );
  AO22X1 U3468 ( .IN1(n6978), .IN2(n6448), .IN3(\FIFO[78][10] ), .IN4(n6450), 
        .Q(n2045) );
  AO22X1 U3469 ( .IN1(n6967), .IN2(n6448), .IN3(\FIFO[78][11] ), .IN4(n6450), 
        .Q(n2046) );
  AO22X1 U3470 ( .IN1(n6956), .IN2(n6448), .IN3(\FIFO[78][12] ), .IN4(n6451), 
        .Q(n2047) );
  AO22X1 U3471 ( .IN1(n6945), .IN2(n6448), .IN3(\FIFO[78][13] ), .IN4(n6451), 
        .Q(n2048) );
  AO22X1 U3472 ( .IN1(n6934), .IN2(n6447), .IN3(\FIFO[78][14] ), .IN4(n6451), 
        .Q(n2049) );
  AO22X1 U3473 ( .IN1(n6923), .IN2(n6447), .IN3(\FIFO[78][15] ), .IN4(n6451), 
        .Q(n2050) );
  AO22X1 U3474 ( .IN1(n6912), .IN2(n6447), .IN3(\FIFO[78][16] ), .IN4(n6451), 
        .Q(n2051) );
  AO22X1 U3475 ( .IN1(n6901), .IN2(n6447), .IN3(\FIFO[78][17] ), .IN4(n6451), 
        .Q(n2052) );
  AO22X1 U3476 ( .IN1(n6890), .IN2(n6447), .IN3(\FIFO[78][18] ), .IN4(n6451), 
        .Q(n2053) );
  AO22X1 U3477 ( .IN1(n6879), .IN2(n6447), .IN3(\FIFO[78][19] ), .IN4(n6451), 
        .Q(n2054) );
  AO22X1 U3478 ( .IN1(n6868), .IN2(n6447), .IN3(\FIFO[78][20] ), .IN4(n6451), 
        .Q(n2055) );
  AO22X1 U3479 ( .IN1(n6857), .IN2(n6449), .IN3(\FIFO[78][21] ), .IN4(n6451), 
        .Q(n2056) );
  AO22X1 U3483 ( .IN1(n6846), .IN2(n6448), .IN3(\FIFO[78][22] ), .IN4(n6451), 
        .Q(n2057) );
  AO22X1 U3489 ( .IN1(n6835), .IN2(n6447), .IN3(\FIFO[78][23] ), .IN4(n6451), 
        .Q(n2058) );
  AO22X1 U3490 ( .IN1(n7094), .IN2(n6431), .IN3(\FIFO[75][0] ), .IN4(n6432), 
        .Q(n2131) );
  AO22X1 U3491 ( .IN1(n7077), .IN2(n6431), .IN3(\FIFO[75][1] ), .IN4(n6432), 
        .Q(n2132) );
  AO22X1 U3492 ( .IN1(n7066), .IN2(n6431), .IN3(\FIFO[75][2] ), .IN4(n6432), 
        .Q(n2133) );
  AO22X1 U3493 ( .IN1(n7055), .IN2(n6431), .IN3(\FIFO[75][3] ), .IN4(n6432), 
        .Q(n2134) );
  AO22X1 U3494 ( .IN1(n7044), .IN2(n6431), .IN3(\FIFO[75][4] ), .IN4(n6432), 
        .Q(n2135) );
  AO22X1 U3495 ( .IN1(n7033), .IN2(n6431), .IN3(\FIFO[75][5] ), .IN4(n6432), 
        .Q(n2136) );
  AO22X1 U3496 ( .IN1(n7022), .IN2(n6431), .IN3(\FIFO[75][6] ), .IN4(n6432), 
        .Q(n2137) );
  AO22X1 U3497 ( .IN1(n7011), .IN2(n6430), .IN3(\FIFO[75][7] ), .IN4(n6432), 
        .Q(n2138) );
  AO22X1 U3498 ( .IN1(n7000), .IN2(n6430), .IN3(\FIFO[75][8] ), .IN4(n6432), 
        .Q(n2139) );
  AO22X1 U3499 ( .IN1(n6989), .IN2(n6430), .IN3(\FIFO[75][9] ), .IN4(n6432), 
        .Q(n2140) );
  AO22X1 U3500 ( .IN1(n6978), .IN2(n6430), .IN3(\FIFO[75][10] ), .IN4(n6432), 
        .Q(n2141) );
  AO22X1 U3501 ( .IN1(n6967), .IN2(n6430), .IN3(\FIFO[75][11] ), .IN4(n6432), 
        .Q(n2142) );
  AO22X1 U3502 ( .IN1(n6956), .IN2(n6430), .IN3(\FIFO[75][12] ), .IN4(n6433), 
        .Q(n2143) );
  AO22X1 U3503 ( .IN1(n6945), .IN2(n6430), .IN3(\FIFO[75][13] ), .IN4(n6433), 
        .Q(n2144) );
  AO22X1 U3504 ( .IN1(n6934), .IN2(n6429), .IN3(\FIFO[75][14] ), .IN4(n6433), 
        .Q(n2145) );
  AO22X1 U3505 ( .IN1(n6923), .IN2(n6429), .IN3(\FIFO[75][15] ), .IN4(n6433), 
        .Q(n2146) );
  AO22X1 U3506 ( .IN1(n6912), .IN2(n6429), .IN3(\FIFO[75][16] ), .IN4(n6433), 
        .Q(n2147) );
  AO22X1 U3507 ( .IN1(n6901), .IN2(n6429), .IN3(\FIFO[75][17] ), .IN4(n6433), 
        .Q(n2148) );
  AO22X1 U3508 ( .IN1(n6890), .IN2(n6429), .IN3(\FIFO[75][18] ), .IN4(n6433), 
        .Q(n2149) );
  AO22X1 U3509 ( .IN1(n6879), .IN2(n6429), .IN3(\FIFO[75][19] ), .IN4(n6433), 
        .Q(n2150) );
  AO22X1 U3510 ( .IN1(n6868), .IN2(n6429), .IN3(\FIFO[75][20] ), .IN4(n6433), 
        .Q(n2151) );
  AO22X1 U3511 ( .IN1(n6857), .IN2(n6431), .IN3(\FIFO[75][21] ), .IN4(n6433), 
        .Q(n2152) );
  AO22X1 U3512 ( .IN1(n6846), .IN2(n6430), .IN3(\FIFO[75][22] ), .IN4(n6433), 
        .Q(n2153) );
  AO22X1 U3524 ( .IN1(n6835), .IN2(n6429), .IN3(\FIFO[75][23] ), .IN4(n6433), 
        .Q(n2154) );
  AO22X1 U3558 ( .IN1(n7094), .IN2(n6425), .IN3(\FIFO[74][0] ), .IN4(n6426), 
        .Q(n2163) );
  AO22X1 U3567 ( .IN1(n7077), .IN2(n6425), .IN3(\FIFO[74][1] ), .IN4(n6426), 
        .Q(n2164) );
  AO22X1 U3588 ( .IN1(n7066), .IN2(n6425), .IN3(\FIFO[74][2] ), .IN4(n6426), 
        .Q(n2165) );
  AO22X1 U3589 ( .IN1(n7055), .IN2(n6425), .IN3(\FIFO[74][3] ), .IN4(n6426), 
        .Q(n2166) );
  AO22X1 U3590 ( .IN1(n7044), .IN2(n6425), .IN3(\FIFO[74][4] ), .IN4(n6426), 
        .Q(n2167) );
  AO22X1 U3591 ( .IN1(n7033), .IN2(n6425), .IN3(\FIFO[74][5] ), .IN4(n6426), 
        .Q(n2168) );
  AO22X1 U3592 ( .IN1(n7022), .IN2(n6425), .IN3(\FIFO[74][6] ), .IN4(n6426), 
        .Q(n2169) );
  AO22X1 U3593 ( .IN1(n7011), .IN2(n6424), .IN3(\FIFO[74][7] ), .IN4(n6426), 
        .Q(n2170) );
  AO22X1 U3594 ( .IN1(n7000), .IN2(n6424), .IN3(\FIFO[74][8] ), .IN4(n6426), 
        .Q(n2171) );
  AO22X1 U3595 ( .IN1(n6989), .IN2(n6424), .IN3(\FIFO[74][9] ), .IN4(n6426), 
        .Q(n2172) );
  AO22X1 U3596 ( .IN1(n6978), .IN2(n6424), .IN3(\FIFO[74][10] ), .IN4(n6426), 
        .Q(n2173) );
  AO22X1 U3597 ( .IN1(n6967), .IN2(n6424), .IN3(\FIFO[74][11] ), .IN4(n6426), 
        .Q(n2174) );
  AO22X1 U3598 ( .IN1(n6956), .IN2(n6424), .IN3(\FIFO[74][12] ), .IN4(n6427), 
        .Q(n2175) );
  AO22X1 U3599 ( .IN1(n6945), .IN2(n6424), .IN3(\FIFO[74][13] ), .IN4(n6427), 
        .Q(n2176) );
  AO22X1 U3600 ( .IN1(n6934), .IN2(n6423), .IN3(\FIFO[74][14] ), .IN4(n6427), 
        .Q(n2177) );
  AO22X1 U3601 ( .IN1(n6923), .IN2(n6423), .IN3(\FIFO[74][15] ), .IN4(n6427), 
        .Q(n2178) );
  AO22X1 U3602 ( .IN1(n6912), .IN2(n6423), .IN3(\FIFO[74][16] ), .IN4(n6427), 
        .Q(n2179) );
  AO22X1 U3603 ( .IN1(n6901), .IN2(n6423), .IN3(\FIFO[74][17] ), .IN4(n6427), 
        .Q(n2180) );
  AO22X1 U3604 ( .IN1(n6890), .IN2(n6423), .IN3(\FIFO[74][18] ), .IN4(n6427), 
        .Q(n2181) );
  AO22X1 U3605 ( .IN1(n6879), .IN2(n6423), .IN3(\FIFO[74][19] ), .IN4(n6427), 
        .Q(n2182) );
  AO22X1 U3606 ( .IN1(n6868), .IN2(n6423), .IN3(\FIFO[74][20] ), .IN4(n6427), 
        .Q(n2183) );
  AO22X1 U3607 ( .IN1(n6857), .IN2(n6425), .IN3(\FIFO[74][21] ), .IN4(n6427), 
        .Q(n2184) );
  AO22X1 U3608 ( .IN1(n6846), .IN2(n6424), .IN3(\FIFO[74][22] ), .IN4(n6427), 
        .Q(n2185) );
  AO22X1 U3609 ( .IN1(n6835), .IN2(n6423), .IN3(\FIFO[74][23] ), .IN4(n6427), 
        .Q(n2186) );
  AO22X1 U3610 ( .IN1(n7093), .IN2(n6407), .IN3(\FIFO[71][0] ), .IN4(n6408), 
        .Q(n2259) );
  AO22X1 U3611 ( .IN1(n7076), .IN2(n6406), .IN3(\FIFO[71][1] ), .IN4(n6408), 
        .Q(n2260) );
  AO22X1 U3616 ( .IN1(n7065), .IN2(n6405), .IN3(\FIFO[71][2] ), .IN4(n6408), 
        .Q(n2261) );
  AO22X1 U3621 ( .IN1(n7054), .IN2(n6407), .IN3(\FIFO[71][3] ), .IN4(n6408), 
        .Q(n2262) );
  AO22X1 U3622 ( .IN1(n7043), .IN2(n6406), .IN3(\FIFO[71][4] ), .IN4(n6408), 
        .Q(n2263) );
  AO22X1 U3623 ( .IN1(n7032), .IN2(n6405), .IN3(\FIFO[71][5] ), .IN4(n6408), 
        .Q(n2264) );
  AO22X1 U3624 ( .IN1(n7021), .IN2(n6407), .IN3(\FIFO[71][6] ), .IN4(n6408), 
        .Q(n2265) );
  AO22X1 U3625 ( .IN1(n7010), .IN2(n6407), .IN3(\FIFO[71][7] ), .IN4(n6408), 
        .Q(n2266) );
  AO22X1 U3626 ( .IN1(n6999), .IN2(n6407), .IN3(\FIFO[71][8] ), .IN4(n6408), 
        .Q(n2267) );
  AO22X1 U3627 ( .IN1(n6988), .IN2(n6407), .IN3(\FIFO[71][9] ), .IN4(n6408), 
        .Q(n2268) );
  AO22X1 U3628 ( .IN1(n6966), .IN2(n6407), .IN3(\FIFO[71][11] ), .IN4(n6408), 
        .Q(n2270) );
  AO22X1 U3629 ( .IN1(n6955), .IN2(n6407), .IN3(\FIFO[71][12] ), .IN4(n6409), 
        .Q(n2271) );
  AO22X1 U3630 ( .IN1(n6944), .IN2(n6407), .IN3(\FIFO[71][13] ), .IN4(n6409), 
        .Q(n2272) );
  AO22X1 U3631 ( .IN1(n6933), .IN2(n6406), .IN3(\FIFO[71][14] ), .IN4(n6409), 
        .Q(n2273) );
  AO22X1 U3632 ( .IN1(n6922), .IN2(n6406), .IN3(\FIFO[71][15] ), .IN4(n6409), 
        .Q(n2274) );
  AO22X1 U3633 ( .IN1(n6911), .IN2(n6406), .IN3(\FIFO[71][16] ), .IN4(n6409), 
        .Q(n2275) );
  AO22X1 U3634 ( .IN1(n6900), .IN2(n6406), .IN3(\FIFO[71][17] ), .IN4(n6409), 
        .Q(n2276) );
  AO22X1 U3635 ( .IN1(n6889), .IN2(n6406), .IN3(\FIFO[71][18] ), .IN4(n6409), 
        .Q(n2277) );
  AO22X1 U3636 ( .IN1(n6878), .IN2(n6406), .IN3(\FIFO[71][19] ), .IN4(n6409), 
        .Q(n2278) );
  AO22X1 U3637 ( .IN1(n6867), .IN2(n6406), .IN3(\FIFO[71][20] ), .IN4(n6409), 
        .Q(n2279) );
  AO22X1 U3638 ( .IN1(n6856), .IN2(n6405), .IN3(\FIFO[71][21] ), .IN4(n6409), 
        .Q(n2280) );
  AO22X1 U3639 ( .IN1(n6845), .IN2(n6405), .IN3(\FIFO[71][22] ), .IN4(n6409), 
        .Q(n2281) );
  AO22X1 U3640 ( .IN1(n7093), .IN2(n6401), .IN3(\FIFO[70][0] ), .IN4(n6402), 
        .Q(n2291) );
  AO22X1 U3641 ( .IN1(n7076), .IN2(n6401), .IN3(\FIFO[70][1] ), .IN4(n6402), 
        .Q(n2292) );
  AO22X1 U3642 ( .IN1(n7065), .IN2(n6401), .IN3(\FIFO[70][2] ), .IN4(n6402), 
        .Q(n2293) );
  AO22X1 U3643 ( .IN1(n7054), .IN2(n6401), .IN3(\FIFO[70][3] ), .IN4(n6402), 
        .Q(n2294) );
  AO22X1 U3644 ( .IN1(n7043), .IN2(n6401), .IN3(\FIFO[70][4] ), .IN4(n6402), 
        .Q(n2295) );
  AO22X1 U3650 ( .IN1(n7032), .IN2(n6401), .IN3(\FIFO[70][5] ), .IN4(n6402), 
        .Q(n2296) );
  AO22X1 U3660 ( .IN1(n7021), .IN2(n6401), .IN3(\FIFO[70][6] ), .IN4(n6402), 
        .Q(n2297) );
  AO22X1 U3667 ( .IN1(n7010), .IN2(n6400), .IN3(\FIFO[70][7] ), .IN4(n6402), 
        .Q(n2298) );
  AO22X1 U3694 ( .IN1(n6999), .IN2(n6400), .IN3(\FIFO[70][8] ), .IN4(n6402), 
        .Q(n2299) );
  AO22X1 U3720 ( .IN1(n6988), .IN2(n6400), .IN3(\FIFO[70][9] ), .IN4(n6402), 
        .Q(n2300) );
  AO22X1 U3721 ( .IN1(n6977), .IN2(n6400), .IN3(\FIFO[70][10] ), .IN4(n6402), 
        .Q(n2301) );
  AO22X1 U3722 ( .IN1(n6966), .IN2(n6400), .IN3(\FIFO[70][11] ), .IN4(n6402), 
        .Q(n2302) );
  AO22X1 U3723 ( .IN1(n6955), .IN2(n6400), .IN3(\FIFO[70][12] ), .IN4(n6403), 
        .Q(n2303) );
  AO22X1 U3724 ( .IN1(n6944), .IN2(n6400), .IN3(\FIFO[70][13] ), .IN4(n6403), 
        .Q(n2304) );
  AO22X1 U3725 ( .IN1(n6933), .IN2(n6399), .IN3(\FIFO[70][14] ), .IN4(n6403), 
        .Q(n2305) );
  AO22X1 U3726 ( .IN1(n6922), .IN2(n6399), .IN3(\FIFO[70][15] ), .IN4(n6403), 
        .Q(n2306) );
  AO22X1 U3727 ( .IN1(n6911), .IN2(n6399), .IN3(\FIFO[70][16] ), .IN4(n6403), 
        .Q(n2307) );
  AO22X1 U3728 ( .IN1(n6900), .IN2(n6399), .IN3(\FIFO[70][17] ), .IN4(n6403), 
        .Q(n2308) );
  AO22X1 U3729 ( .IN1(n6889), .IN2(n6399), .IN3(\FIFO[70][18] ), .IN4(n6403), 
        .Q(n2309) );
  AO22X1 U3730 ( .IN1(n6878), .IN2(n6399), .IN3(\FIFO[70][19] ), .IN4(n6403), 
        .Q(n2310) );
  AO22X1 U3731 ( .IN1(n6867), .IN2(n6399), .IN3(\FIFO[70][20] ), .IN4(n6403), 
        .Q(n2311) );
  AO22X1 U3732 ( .IN1(n6856), .IN2(n6401), .IN3(\FIFO[70][21] ), .IN4(n6403), 
        .Q(n2312) );
  AO22X1 U3733 ( .IN1(n6845), .IN2(n6400), .IN3(\FIFO[70][22] ), .IN4(n6403), 
        .Q(n2313) );
  AO22X1 U3734 ( .IN1(n6834), .IN2(n6399), .IN3(\FIFO[70][23] ), .IN4(n6403), 
        .Q(n2314) );
  AO22X1 U3735 ( .IN1(n7093), .IN2(n6383), .IN3(\FIFO[67][0] ), .IN4(n6384), 
        .Q(n2387) );
  AO22X1 U3736 ( .IN1(n7076), .IN2(n6383), .IN3(\FIFO[67][1] ), .IN4(n6384), 
        .Q(n2388) );
  AO22X1 U3737 ( .IN1(n7065), .IN2(n6383), .IN3(\FIFO[67][2] ), .IN4(n6384), 
        .Q(n2389) );
  AO22X1 U3738 ( .IN1(n7054), .IN2(n6383), .IN3(\FIFO[67][3] ), .IN4(n6384), 
        .Q(n2390) );
  AO22X1 U3739 ( .IN1(n7043), .IN2(n6383), .IN3(\FIFO[67][4] ), .IN4(n6384), 
        .Q(n2391) );
  AO22X1 U3740 ( .IN1(n7032), .IN2(n6383), .IN3(\FIFO[67][5] ), .IN4(n6384), 
        .Q(n2392) );
  AO22X1 U3741 ( .IN1(n7021), .IN2(n6383), .IN3(\FIFO[67][6] ), .IN4(n6384), 
        .Q(n2393) );
  AO22X1 U3742 ( .IN1(n7010), .IN2(n6382), .IN3(\FIFO[67][7] ), .IN4(n6384), 
        .Q(n2394) );
  AO22X1 U3743 ( .IN1(n6999), .IN2(n6382), .IN3(\FIFO[67][8] ), .IN4(n6384), 
        .Q(n2395) );
  AO22X1 U3753 ( .IN1(n6988), .IN2(n6382), .IN3(\FIFO[67][9] ), .IN4(n6384), 
        .Q(n2396) );
  AO22X1 U3754 ( .IN1(n6977), .IN2(n6382), .IN3(\FIFO[67][10] ), .IN4(n6384), 
        .Q(n2397) );
  AO22X1 U3755 ( .IN1(n6966), .IN2(n6382), .IN3(\FIFO[67][11] ), .IN4(n6384), 
        .Q(n2398) );
  AO22X1 U3756 ( .IN1(n6944), .IN2(n6382), .IN3(\FIFO[67][13] ), .IN4(n6385), 
        .Q(n2400) );
  AO22X1 U3757 ( .IN1(n6933), .IN2(n6383), .IN3(\FIFO[67][14] ), .IN4(n6385), 
        .Q(n2401) );
  AO22X1 U3758 ( .IN1(n6922), .IN2(n6382), .IN3(\FIFO[67][15] ), .IN4(n6385), 
        .Q(n2402) );
  AO22X1 U3759 ( .IN1(n6911), .IN2(n6381), .IN3(\FIFO[67][16] ), .IN4(n6385), 
        .Q(n2403) );
  AO22X1 U3760 ( .IN1(n6900), .IN2(n6383), .IN3(\FIFO[67][17] ), .IN4(n6385), 
        .Q(n2404) );
  AO22X1 U3761 ( .IN1(n6889), .IN2(n6382), .IN3(\FIFO[67][18] ), .IN4(n6385), 
        .Q(n2405) );
  AO22X1 U3762 ( .IN1(n6878), .IN2(n6381), .IN3(\FIFO[67][19] ), .IN4(n6385), 
        .Q(n2406) );
  AO22X1 U3763 ( .IN1(n6867), .IN2(n6383), .IN3(\FIFO[67][20] ), .IN4(n6385), 
        .Q(n2407) );
  AO22X1 U3764 ( .IN1(n6856), .IN2(n6381), .IN3(\FIFO[67][21] ), .IN4(n6385), 
        .Q(n2408) );
  AO22X1 U3765 ( .IN1(n6845), .IN2(n6381), .IN3(\FIFO[67][22] ), .IN4(n6385), 
        .Q(n2409) );
  AO22X1 U3766 ( .IN1(n6834), .IN2(n6381), .IN3(\FIFO[67][23] ), .IN4(n6385), 
        .Q(n2410) );
  AO22X1 U3767 ( .IN1(n7093), .IN2(n6377), .IN3(\FIFO[66][0] ), .IN4(n6378), 
        .Q(n2419) );
  AO22X1 U3768 ( .IN1(n7076), .IN2(n6376), .IN3(\FIFO[66][1] ), .IN4(n6378), 
        .Q(n2420) );
  AO22X1 U3769 ( .IN1(n7065), .IN2(n6375), .IN3(\FIFO[66][2] ), .IN4(n6378), 
        .Q(n2421) );
  AO22X1 U3770 ( .IN1(n7054), .IN2(n6377), .IN3(\FIFO[66][3] ), .IN4(n6378), 
        .Q(n2422) );
  AO22X1 U3771 ( .IN1(n7032), .IN2(n6375), .IN3(\FIFO[66][5] ), .IN4(n6378), 
        .Q(n2424) );
  AO22X1 U3772 ( .IN1(n7021), .IN2(n6377), .IN3(\FIFO[66][6] ), .IN4(n6378), 
        .Q(n2425) );
  AO22X1 U3773 ( .IN1(n7010), .IN2(n6377), .IN3(\FIFO[66][7] ), .IN4(n6378), 
        .Q(n2426) );
  AO22X1 U3774 ( .IN1(n6999), .IN2(n6377), .IN3(\FIFO[66][8] ), .IN4(n6378), 
        .Q(n2427) );
  AO22X1 U3775 ( .IN1(n6988), .IN2(n6377), .IN3(\FIFO[66][9] ), .IN4(n6378), 
        .Q(n2428) );
  AO22X1 U3776 ( .IN1(n6977), .IN2(n6377), .IN3(\FIFO[66][10] ), .IN4(n6378), 
        .Q(n2429) );
  AO22X1 U3783 ( .IN1(n6966), .IN2(n6377), .IN3(\FIFO[66][11] ), .IN4(n6378), 
        .Q(n2430) );
  AO22X1 U3796 ( .IN1(n6955), .IN2(n6377), .IN3(\FIFO[66][12] ), .IN4(n6379), 
        .Q(n2431) );
  AO22X1 U3809 ( .IN1(n6933), .IN2(n6376), .IN3(\FIFO[66][14] ), .IN4(n6379), 
        .Q(n2433) );
  AO22X1 U3817 ( .IN1(n6922), .IN2(n6376), .IN3(\FIFO[66][15] ), .IN4(n6379), 
        .Q(n2434) );
  AO22X1 U3830 ( .IN1(n6911), .IN2(n6376), .IN3(\FIFO[66][16] ), .IN4(n6379), 
        .Q(n2435) );
  AO22X1 U3852 ( .IN1(n6900), .IN2(n6376), .IN3(\FIFO[66][17] ), .IN4(n6379), 
        .Q(n2436) );
  AO22X1 U3853 ( .IN1(n6889), .IN2(n6376), .IN3(\FIFO[66][18] ), .IN4(n6379), 
        .Q(n2437) );
  AO22X1 U3854 ( .IN1(n6878), .IN2(n6376), .IN3(\FIFO[66][19] ), .IN4(n6379), 
        .Q(n2438) );
  AO22X1 U3855 ( .IN1(n6867), .IN2(n6376), .IN3(\FIFO[66][20] ), .IN4(n6379), 
        .Q(n2439) );
  AO22X1 U3856 ( .IN1(n6856), .IN2(n6375), .IN3(\FIFO[66][21] ), .IN4(n6379), 
        .Q(n2440) );
  AO22X1 U3857 ( .IN1(n6845), .IN2(n6375), .IN3(\FIFO[66][22] ), .IN4(n6379), 
        .Q(n2441) );
  AO22X1 U3858 ( .IN1(n6834), .IN2(n6375), .IN3(\FIFO[66][23] ), .IN4(n6379), 
        .Q(n2442) );
  AO22X1 U3859 ( .IN1(n7093), .IN2(n6359), .IN3(\FIFO[63][0] ), .IN4(n6360), 
        .Q(n2515) );
  AO22X1 U3860 ( .IN1(n7076), .IN2(n6359), .IN3(\FIFO[63][1] ), .IN4(n6360), 
        .Q(n2516) );
  AO22X1 U3861 ( .IN1(n7065), .IN2(n6359), .IN3(\FIFO[63][2] ), .IN4(n6360), 
        .Q(n2517) );
  AO22X1 U3862 ( .IN1(n7054), .IN2(n6359), .IN3(\FIFO[63][3] ), .IN4(n6360), 
        .Q(n2518) );
  AO22X1 U3863 ( .IN1(n7043), .IN2(n6359), .IN3(\FIFO[63][4] ), .IN4(n6360), 
        .Q(n2519) );
  AO22X1 U3864 ( .IN1(n7032), .IN2(n6359), .IN3(\FIFO[63][5] ), .IN4(n6360), 
        .Q(n2520) );
  AO22X1 U3865 ( .IN1(n7021), .IN2(n6359), .IN3(\FIFO[63][6] ), .IN4(n6360), 
        .Q(n2521) );
  AO22X1 U3866 ( .IN1(n7010), .IN2(n6358), .IN3(\FIFO[63][7] ), .IN4(n6360), 
        .Q(n2522) );
  AO22X1 U3867 ( .IN1(n6999), .IN2(n6358), .IN3(\FIFO[63][8] ), .IN4(n6360), 
        .Q(n2523) );
  AO22X1 U3868 ( .IN1(n6977), .IN2(n6358), .IN3(\FIFO[63][10] ), .IN4(n6360), 
        .Q(n2525) );
  AO22X1 U3869 ( .IN1(n6966), .IN2(n6358), .IN3(\FIFO[63][11] ), .IN4(n6360), 
        .Q(n2526) );
  AO22X1 U3870 ( .IN1(n6955), .IN2(n6358), .IN3(\FIFO[63][12] ), .IN4(n6361), 
        .Q(n2527) );
  AO22X1 U3871 ( .IN1(n6944), .IN2(n6358), .IN3(\FIFO[63][13] ), .IN4(n6361), 
        .Q(n2528) );
  AO22X1 U3872 ( .IN1(n6922), .IN2(n6358), .IN3(\FIFO[63][15] ), .IN4(n6361), 
        .Q(n2530) );
  AO22X1 U3873 ( .IN1(n6911), .IN2(n6357), .IN3(\FIFO[63][16] ), .IN4(n6361), 
        .Q(n2531) );
  AO22X1 U3874 ( .IN1(n6900), .IN2(n6359), .IN3(\FIFO[63][17] ), .IN4(n6361), 
        .Q(n2532) );
  AO22X1 U3875 ( .IN1(n6889), .IN2(n6358), .IN3(\FIFO[63][18] ), .IN4(n6361), 
        .Q(n2533) );
  AO22X1 U3885 ( .IN1(n6878), .IN2(n6357), .IN3(\FIFO[63][19] ), .IN4(n6361), 
        .Q(n2534) );
  AO22X1 U3886 ( .IN1(n6867), .IN2(n6359), .IN3(\FIFO[63][20] ), .IN4(n6361), 
        .Q(n2535) );
  AO22X1 U3887 ( .IN1(n6856), .IN2(n6357), .IN3(\FIFO[63][21] ), .IN4(n6361), 
        .Q(n2536) );
  AO22X1 U3888 ( .IN1(n6845), .IN2(n6357), .IN3(\FIFO[63][22] ), .IN4(n6361), 
        .Q(n2537) );
  AO22X1 U3889 ( .IN1(n6834), .IN2(n6357), .IN3(\FIFO[63][23] ), .IN4(n6361), 
        .Q(n2538) );
  AO22X1 U3890 ( .IN1(n7093), .IN2(n6353), .IN3(\FIFO[62][0] ), .IN4(n6354), 
        .Q(n2547) );
  AO22X1 U3891 ( .IN1(n7076), .IN2(n6352), .IN3(\FIFO[62][1] ), .IN4(n6354), 
        .Q(n2548) );
  AO22X1 U3892 ( .IN1(n7065), .IN2(n6351), .IN3(\FIFO[62][2] ), .IN4(n6354), 
        .Q(n2549) );
  AO22X1 U3893 ( .IN1(n7054), .IN2(n6353), .IN3(\FIFO[62][3] ), .IN4(n6354), 
        .Q(n2550) );
  AO22X1 U3894 ( .IN1(n7043), .IN2(n6352), .IN3(\FIFO[62][4] ), .IN4(n6354), 
        .Q(n2551) );
  AO22X1 U3895 ( .IN1(n7032), .IN2(n6351), .IN3(\FIFO[62][5] ), .IN4(n6354), 
        .Q(n2552) );
  AO22X1 U3896 ( .IN1(n7021), .IN2(n6353), .IN3(\FIFO[62][6] ), .IN4(n6354), 
        .Q(n2553) );
  AO22X1 U3897 ( .IN1(n7010), .IN2(n6353), .IN3(\FIFO[62][7] ), .IN4(n6354), 
        .Q(n2554) );
  AO22X1 U3898 ( .IN1(n6999), .IN2(n6353), .IN3(\FIFO[62][8] ), .IN4(n6354), 
        .Q(n2555) );
  AO22X1 U3899 ( .IN1(n6988), .IN2(n6353), .IN3(\FIFO[62][9] ), .IN4(n6354), 
        .Q(n2556) );
  AO22X1 U3900 ( .IN1(n6977), .IN2(n6353), .IN3(\FIFO[62][10] ), .IN4(n6354), 
        .Q(n2557) );
  AO22X1 U3901 ( .IN1(n6966), .IN2(n6353), .IN3(\FIFO[62][11] ), .IN4(n6354), 
        .Q(n2558) );
  AO22X1 U3902 ( .IN1(n6955), .IN2(n6353), .IN3(\FIFO[62][12] ), .IN4(n6355), 
        .Q(n2559) );
  AO22X1 U3903 ( .IN1(n6944), .IN2(n6353), .IN3(\FIFO[62][13] ), .IN4(n6355), 
        .Q(n2560) );
  AO22X1 U3904 ( .IN1(n6933), .IN2(n6352), .IN3(\FIFO[62][14] ), .IN4(n6355), 
        .Q(n2561) );
  AO22X1 U3905 ( .IN1(n6911), .IN2(n6352), .IN3(\FIFO[62][16] ), .IN4(n6355), 
        .Q(n2563) );
  AO22X1 U3906 ( .IN1(n6900), .IN2(n6352), .IN3(\FIFO[62][17] ), .IN4(n6355), 
        .Q(n2564) );
  AO22X1 U3907 ( .IN1(n6889), .IN2(n6352), .IN3(\FIFO[62][18] ), .IN4(n6355), 
        .Q(n2565) );
  AO22X1 U3908 ( .IN1(n6878), .IN2(n6352), .IN3(\FIFO[62][19] ), .IN4(n6355), 
        .Q(n2566) );
  AO22X1 U3929 ( .IN1(n6867), .IN2(n6352), .IN3(\FIFO[62][20] ), .IN4(n6355), 
        .Q(n2567) );
  AO22X1 U3934 ( .IN1(n6856), .IN2(n6351), .IN3(\FIFO[62][21] ), .IN4(n6355), 
        .Q(n2568) );
  AO22X1 U3942 ( .IN1(n6845), .IN2(n6351), .IN3(\FIFO[62][22] ), .IN4(n6355), 
        .Q(n2569) );
  AO22X1 U3956 ( .IN1(n6834), .IN2(n6351), .IN3(\FIFO[62][23] ), .IN4(n6355), 
        .Q(n2570) );
  AO22X1 U3968 ( .IN1(n7092), .IN2(n6335), .IN3(\FIFO[59][0] ), .IN4(n6336), 
        .Q(n2643) );
  AO22X1 U3976 ( .IN1(n7075), .IN2(n6335), .IN3(\FIFO[59][1] ), .IN4(n6336), 
        .Q(n2644) );
  AO22X1 U3984 ( .IN1(n7064), .IN2(n6335), .IN3(\FIFO[59][2] ), .IN4(n6336), 
        .Q(n2645) );
  AO22X1 U3985 ( .IN1(n7053), .IN2(n6335), .IN3(\FIFO[59][3] ), .IN4(n6336), 
        .Q(n2646) );
  AO22X1 U3986 ( .IN1(n7042), .IN2(n6335), .IN3(\FIFO[59][4] ), .IN4(n6336), 
        .Q(n2647) );
  AO22X1 U3987 ( .IN1(n7031), .IN2(n6335), .IN3(\FIFO[59][5] ), .IN4(n6336), 
        .Q(n2648) );
  AO22X1 U3988 ( .IN1(n7020), .IN2(n6335), .IN3(\FIFO[59][6] ), .IN4(n6336), 
        .Q(n2649) );
  AO22X1 U3989 ( .IN1(n7009), .IN2(n6334), .IN3(\FIFO[59][7] ), .IN4(n6336), 
        .Q(n2650) );
  AO22X1 U3990 ( .IN1(n6998), .IN2(n6334), .IN3(\FIFO[59][8] ), .IN4(n6336), 
        .Q(n2651) );
  AO22X1 U3991 ( .IN1(n6987), .IN2(n6334), .IN3(\FIFO[59][9] ), .IN4(n6336), 
        .Q(n2652) );
  AO22X1 U3992 ( .IN1(n6976), .IN2(n6334), .IN3(\FIFO[59][10] ), .IN4(n6336), 
        .Q(n2653) );
  AO22X1 U3993 ( .IN1(n6965), .IN2(n6334), .IN3(\FIFO[59][11] ), .IN4(n6336), 
        .Q(n2654) );
  AO22X1 U3994 ( .IN1(n6954), .IN2(n6334), .IN3(\FIFO[59][12] ), .IN4(n6337), 
        .Q(n2655) );
  AO22X1 U3995 ( .IN1(n6943), .IN2(n6334), .IN3(\FIFO[59][13] ), .IN4(n6337), 
        .Q(n2656) );
  AO22X1 U3996 ( .IN1(n6932), .IN2(n6333), .IN3(\FIFO[59][14] ), .IN4(n6337), 
        .Q(n2657) );
  AO22X1 U3997 ( .IN1(n6921), .IN2(n6333), .IN3(\FIFO[59][15] ), .IN4(n6337), 
        .Q(n2658) );
  AO22X1 U3998 ( .IN1(n6910), .IN2(n6333), .IN3(\FIFO[59][16] ), .IN4(n6337), 
        .Q(n2659) );
  AO22X1 U3999 ( .IN1(n6899), .IN2(n6333), .IN3(\FIFO[59][17] ), .IN4(n6337), 
        .Q(n2660) );
  AO22X1 U4000 ( .IN1(n6888), .IN2(n6333), .IN3(\FIFO[59][18] ), .IN4(n6337), 
        .Q(n2661) );
  AO22X1 U4001 ( .IN1(n6877), .IN2(n6333), .IN3(\FIFO[59][19] ), .IN4(n6337), 
        .Q(n2662) );
  AO22X1 U4002 ( .IN1(n6866), .IN2(n6333), .IN3(\FIFO[59][20] ), .IN4(n6337), 
        .Q(n2663) );
  AO22X1 U4003 ( .IN1(n6855), .IN2(n6335), .IN3(\FIFO[59][21] ), .IN4(n6337), 
        .Q(n2664) );
  AO22X1 U4004 ( .IN1(n6844), .IN2(n6334), .IN3(\FIFO[59][22] ), .IN4(n6337), 
        .Q(n2665) );
  AO22X1 U4005 ( .IN1(n6833), .IN2(n6333), .IN3(\FIFO[59][23] ), .IN4(n6337), 
        .Q(n2666) );
  AO22X1 U4006 ( .IN1(n7092), .IN2(n6329), .IN3(\FIFO[58][0] ), .IN4(n6330), 
        .Q(n2675) );
  AO22X1 U4007 ( .IN1(n7075), .IN2(n6329), .IN3(\FIFO[58][1] ), .IN4(n6330), 
        .Q(n2676) );
  AO22X1 U4008 ( .IN1(n7064), .IN2(n6329), .IN3(\FIFO[58][2] ), .IN4(n6330), 
        .Q(n2677) );
  AO22X1 U4017 ( .IN1(n7053), .IN2(n6329), .IN3(\FIFO[58][3] ), .IN4(n6330), 
        .Q(n2678) );
  AO22X1 U4018 ( .IN1(n7042), .IN2(n6329), .IN3(\FIFO[58][4] ), .IN4(n6330), 
        .Q(n2679) );
  AO22X1 U4019 ( .IN1(n7031), .IN2(n6329), .IN3(\FIFO[58][5] ), .IN4(n6330), 
        .Q(n2680) );
  AO22X1 U4020 ( .IN1(n7020), .IN2(n6329), .IN3(\FIFO[58][6] ), .IN4(n6330), 
        .Q(n2681) );
  AO22X1 U4021 ( .IN1(n7009), .IN2(n6328), .IN3(\FIFO[58][7] ), .IN4(n6330), 
        .Q(n2682) );
  AO22X1 U4022 ( .IN1(n6998), .IN2(n6328), .IN3(\FIFO[58][8] ), .IN4(n6330), 
        .Q(n2683) );
  AO22X1 U4023 ( .IN1(n6987), .IN2(n6328), .IN3(\FIFO[58][9] ), .IN4(n6330), 
        .Q(n2684) );
  AO22X1 U4024 ( .IN1(n6965), .IN2(n6328), .IN3(\FIFO[58][11] ), .IN4(n6330), 
        .Q(n2686) );
  AO22X1 U4025 ( .IN1(n6954), .IN2(n6328), .IN3(\FIFO[58][12] ), .IN4(n6331), 
        .Q(n2687) );
  AO22X1 U4026 ( .IN1(n6943), .IN2(n6328), .IN3(\FIFO[58][13] ), .IN4(n6331), 
        .Q(n2688) );
  AO22X1 U4027 ( .IN1(n6932), .IN2(n6329), .IN3(\FIFO[58][14] ), .IN4(n6331), 
        .Q(n2689) );
  AO22X1 U4028 ( .IN1(n6921), .IN2(n6328), .IN3(\FIFO[58][15] ), .IN4(n6331), 
        .Q(n2690) );
  AO22X1 U4029 ( .IN1(n6899), .IN2(n6329), .IN3(\FIFO[58][17] ), .IN4(n6331), 
        .Q(n2692) );
  AO22X1 U4030 ( .IN1(n6888), .IN2(n6328), .IN3(\FIFO[58][18] ), .IN4(n6331), 
        .Q(n2693) );
  AO22X1 U4031 ( .IN1(n6877), .IN2(n6327), .IN3(\FIFO[58][19] ), .IN4(n6331), 
        .Q(n2694) );
  AO22X1 U4032 ( .IN1(n6866), .IN2(n6329), .IN3(\FIFO[58][20] ), .IN4(n6331), 
        .Q(n2695) );
  AO22X1 U4033 ( .IN1(n6855), .IN2(n6327), .IN3(\FIFO[58][21] ), .IN4(n6331), 
        .Q(n2696) );
  AO22X1 U4034 ( .IN1(n6844), .IN2(n6327), .IN3(\FIFO[58][22] ), .IN4(n6331), 
        .Q(n2697) );
  AO22X1 U4035 ( .IN1(n6833), .IN2(n6327), .IN3(\FIFO[58][23] ), .IN4(n6331), 
        .Q(n2698) );
  AO22X1 U4036 ( .IN1(n7092), .IN2(n6311), .IN3(\FIFO[55][0] ), .IN4(n6312), 
        .Q(n2771) );
  AO22X1 U4037 ( .IN1(n7075), .IN2(n6311), .IN3(\FIFO[55][1] ), .IN4(n6312), 
        .Q(n2772) );
  AO22X1 U4038 ( .IN1(n7064), .IN2(n6311), .IN3(\FIFO[55][2] ), .IN4(n6312), 
        .Q(n2773) );
  AO22X1 U4039 ( .IN1(n7053), .IN2(n6311), .IN3(\FIFO[55][3] ), .IN4(n6312), 
        .Q(n2774) );
  AO22X1 U4040 ( .IN1(n7042), .IN2(n6311), .IN3(\FIFO[55][4] ), .IN4(n6312), 
        .Q(n2775) );
  AO22X1 U4041 ( .IN1(n7031), .IN2(n6311), .IN3(\FIFO[55][5] ), .IN4(n6312), 
        .Q(n2776) );
  AO22X1 U4042 ( .IN1(n7020), .IN2(n6311), .IN3(\FIFO[55][6] ), .IN4(n6312), 
        .Q(n2777) );
  AO22X1 U4051 ( .IN1(n7009), .IN2(n6310), .IN3(\FIFO[55][7] ), .IN4(n6312), 
        .Q(n2778) );
  AO22X1 U4052 ( .IN1(n6998), .IN2(n6310), .IN3(\FIFO[55][8] ), .IN4(n6312), 
        .Q(n2779) );
  AO22X1 U4059 ( .IN1(n6987), .IN2(n6310), .IN3(\FIFO[55][9] ), .IN4(n6312), 
        .Q(n2780) );
  AO22X1 U4071 ( .IN1(n6976), .IN2(n6310), .IN3(\FIFO[55][10] ), .IN4(n6312), 
        .Q(n2781) );
  AO22X1 U4079 ( .IN1(n6965), .IN2(n6310), .IN3(\FIFO[55][11] ), .IN4(n6312), 
        .Q(n2782) );
  AO22X1 U4094 ( .IN1(n6954), .IN2(n6310), .IN3(\FIFO[55][12] ), .IN4(n6313), 
        .Q(n2783) );
  AO22X1 U4106 ( .IN1(n6943), .IN2(n6310), .IN3(\FIFO[55][13] ), .IN4(n6313), 
        .Q(n2784) );
  AO22X1 U4114 ( .IN1(n6932), .IN2(n6309), .IN3(\FIFO[55][14] ), .IN4(n6313), 
        .Q(n2785) );
  AO22X1 U4121 ( .IN1(n6921), .IN2(n6309), .IN3(\FIFO[55][15] ), .IN4(n6313), 
        .Q(n2786) );
  AO22X1 U4122 ( .IN1(n6910), .IN2(n6309), .IN3(\FIFO[55][16] ), .IN4(n6313), 
        .Q(n2787) );
  AO22X1 U4123 ( .IN1(n6899), .IN2(n6309), .IN3(\FIFO[55][17] ), .IN4(n6313), 
        .Q(n2788) );
  AO22X1 U4124 ( .IN1(n6888), .IN2(n6309), .IN3(\FIFO[55][18] ), .IN4(n6313), 
        .Q(n2789) );
  AO22X1 U4125 ( .IN1(n6877), .IN2(n6309), .IN3(\FIFO[55][19] ), .IN4(n6313), 
        .Q(n2790) );
  AO22X1 U4126 ( .IN1(n6866), .IN2(n6309), .IN3(\FIFO[55][20] ), .IN4(n6313), 
        .Q(n2791) );
  AO22X1 U4127 ( .IN1(n6855), .IN2(n6311), .IN3(\FIFO[55][21] ), .IN4(n6313), 
        .Q(n2792) );
  AO22X1 U4128 ( .IN1(n6844), .IN2(n6310), .IN3(\FIFO[55][22] ), .IN4(n6313), 
        .Q(n2793) );
  AO22X1 U4129 ( .IN1(n6833), .IN2(n6309), .IN3(\FIFO[55][23] ), .IN4(n6313), 
        .Q(n2794) );
  AO22X1 U4130 ( .IN1(n7092), .IN2(n6305), .IN3(\FIFO[54][0] ), .IN4(n6306), 
        .Q(n2803) );
  AO22X1 U4131 ( .IN1(n7075), .IN2(n6305), .IN3(\FIFO[54][1] ), .IN4(n6306), 
        .Q(n2804) );
  AO22X1 U4132 ( .IN1(n7064), .IN2(n6305), .IN3(\FIFO[54][2] ), .IN4(n6306), 
        .Q(n2805) );
  AO22X1 U4133 ( .IN1(n7053), .IN2(n6305), .IN3(\FIFO[54][3] ), .IN4(n6306), 
        .Q(n2806) );
  AO22X1 U4134 ( .IN1(n7042), .IN2(n6305), .IN3(\FIFO[54][4] ), .IN4(n6306), 
        .Q(n2807) );
  AO22X1 U4135 ( .IN1(n7031), .IN2(n6305), .IN3(\FIFO[54][5] ), .IN4(n6306), 
        .Q(n2808) );
  AO22X1 U4136 ( .IN1(n7020), .IN2(n6305), .IN3(\FIFO[54][6] ), .IN4(n6306), 
        .Q(n2809) );
  AO22X1 U4137 ( .IN1(n7009), .IN2(n6304), .IN3(\FIFO[54][7] ), .IN4(n6306), 
        .Q(n2810) );
  AO22X1 U4138 ( .IN1(n6998), .IN2(n6304), .IN3(\FIFO[54][8] ), .IN4(n6306), 
        .Q(n2811) );
  AO22X1 U4139 ( .IN1(n6987), .IN2(n6304), .IN3(\FIFO[54][9] ), .IN4(n6306), 
        .Q(n2812) );
  AO22X1 U4140 ( .IN1(n6976), .IN2(n6304), .IN3(\FIFO[54][10] ), .IN4(n6306), 
        .Q(n2813) );
  AO22X1 U4141 ( .IN1(n6965), .IN2(n6304), .IN3(\FIFO[54][11] ), .IN4(n6306), 
        .Q(n2814) );
  AO22X1 U4142 ( .IN1(n6954), .IN2(n6304), .IN3(\FIFO[54][12] ), .IN4(n6307), 
        .Q(n2815) );
  AO22X1 U4143 ( .IN1(n6943), .IN2(n6304), .IN3(\FIFO[54][13] ), .IN4(n6307), 
        .Q(n2816) );
  AO22X1 U4144 ( .IN1(n6932), .IN2(n6303), .IN3(\FIFO[54][14] ), .IN4(n6307), 
        .Q(n2817) );
  AO22X1 U4153 ( .IN1(n6921), .IN2(n6303), .IN3(\FIFO[54][15] ), .IN4(n6307), 
        .Q(n2818) );
  AO22X1 U4154 ( .IN1(n6910), .IN2(n6303), .IN3(\FIFO[54][16] ), .IN4(n6307), 
        .Q(n2819) );
  AO22X1 U4155 ( .IN1(n6899), .IN2(n6303), .IN3(\FIFO[54][17] ), .IN4(n6307), 
        .Q(n2820) );
  AO22X1 U4156 ( .IN1(n6888), .IN2(n6303), .IN3(\FIFO[54][18] ), .IN4(n6307), 
        .Q(n2821) );
  AO22X1 U4157 ( .IN1(n6877), .IN2(n6303), .IN3(\FIFO[54][19] ), .IN4(n6307), 
        .Q(n2822) );
  AO22X1 U4158 ( .IN1(n6866), .IN2(n6303), .IN3(\FIFO[54][20] ), .IN4(n6307), 
        .Q(n2823) );
  AO22X1 U4159 ( .IN1(n6855), .IN2(n6305), .IN3(\FIFO[54][21] ), .IN4(n6307), 
        .Q(n2824) );
  AO22X1 U4160 ( .IN1(n6844), .IN2(n6304), .IN3(\FIFO[54][22] ), .IN4(n6307), 
        .Q(n2825) );
  AO22X1 U4161 ( .IN1(n6833), .IN2(n6303), .IN3(\FIFO[54][23] ), .IN4(n6307), 
        .Q(n2826) );
  AO22X1 U4162 ( .IN1(n7092), .IN2(n6287), .IN3(\FIFO[51][0] ), .IN4(n6288), 
        .Q(n2899) );
  AO22X1 U4163 ( .IN1(n7075), .IN2(n6287), .IN3(\FIFO[51][1] ), .IN4(n6288), 
        .Q(n2900) );
  AO22X1 U4164 ( .IN1(n7064), .IN2(n6287), .IN3(\FIFO[51][2] ), .IN4(n6288), 
        .Q(n2901) );
  AO22X1 U4165 ( .IN1(n7053), .IN2(n6287), .IN3(\FIFO[51][3] ), .IN4(n6288), 
        .Q(n2902) );
  AO22X1 U4166 ( .IN1(n7042), .IN2(n6287), .IN3(\FIFO[51][4] ), .IN4(n6288), 
        .Q(n2903) );
  AO22X1 U4167 ( .IN1(n7031), .IN2(n6287), .IN3(\FIFO[51][5] ), .IN4(n6288), 
        .Q(n2904) );
  AO22X1 U4168 ( .IN1(n7020), .IN2(n6287), .IN3(\FIFO[51][6] ), .IN4(n6288), 
        .Q(n2905) );
  AO22X1 U4169 ( .IN1(n7009), .IN2(n6286), .IN3(\FIFO[51][7] ), .IN4(n6288), 
        .Q(n2906) );
  AO22X1 U4170 ( .IN1(n6998), .IN2(n6286), .IN3(\FIFO[51][8] ), .IN4(n6288), 
        .Q(n2907) );
  AO22X1 U4171 ( .IN1(n6987), .IN2(n6286), .IN3(\FIFO[51][9] ), .IN4(n6288), 
        .Q(n2908) );
  AO22X1 U4172 ( .IN1(n6976), .IN2(n6286), .IN3(\FIFO[51][10] ), .IN4(n6288), 
        .Q(n2909) );
  AO22X1 U4173 ( .IN1(n6965), .IN2(n6286), .IN3(\FIFO[51][11] ), .IN4(n6288), 
        .Q(n2910) );
  AO22X1 U4174 ( .IN1(n6954), .IN2(n6286), .IN3(\FIFO[51][12] ), .IN4(n6289), 
        .Q(n2911) );
  AO22X1 U4175 ( .IN1(n6943), .IN2(n6286), .IN3(\FIFO[51][13] ), .IN4(n6289), 
        .Q(n2912) );
  AO22X1 U4176 ( .IN1(n6932), .IN2(n6285), .IN3(\FIFO[51][14] ), .IN4(n6289), 
        .Q(n2913) );
  AO22X1 U4177 ( .IN1(n6921), .IN2(n6285), .IN3(\FIFO[51][15] ), .IN4(n6289), 
        .Q(n2914) );
  AO22X1 U4178 ( .IN1(n6910), .IN2(n6285), .IN3(\FIFO[51][16] ), .IN4(n6289), 
        .Q(n2915) );
  AO22X1 U4187 ( .IN1(n6899), .IN2(n6285), .IN3(\FIFO[51][17] ), .IN4(n6289), 
        .Q(n2916) );
  AO22X1 U4188 ( .IN1(n6888), .IN2(n6285), .IN3(\FIFO[51][18] ), .IN4(n6289), 
        .Q(n2917) );
  AO22X1 U4196 ( .IN1(n6877), .IN2(n6285), .IN3(\FIFO[51][19] ), .IN4(n6289), 
        .Q(n2918) );
  AO22X1 U4207 ( .IN1(n6866), .IN2(n6285), .IN3(\FIFO[51][20] ), .IN4(n6289), 
        .Q(n2919) );
  AO22X1 U4221 ( .IN1(n6855), .IN2(n6287), .IN3(\FIFO[51][21] ), .IN4(n6289), 
        .Q(n2920) );
  AO22X1 U4222 ( .IN1(n6844), .IN2(n6286), .IN3(\FIFO[51][22] ), .IN4(n6289), 
        .Q(n2921) );
  AO22X1 U4236 ( .IN1(n6833), .IN2(n6285), .IN3(\FIFO[51][23] ), .IN4(n6289), 
        .Q(n2922) );
  AO22X1 U4243 ( .IN1(n7092), .IN2(n6281), .IN3(\FIFO[50][0] ), .IN4(n6282), 
        .Q(n2931) );
  AO22X1 U4251 ( .IN1(n7075), .IN2(n6281), .IN3(\FIFO[50][1] ), .IN4(n6282), 
        .Q(n2932) );
  AO22X1 U4257 ( .IN1(n7064), .IN2(n6281), .IN3(\FIFO[50][2] ), .IN4(n6282), 
        .Q(n2933) );
  AO22X1 U4258 ( .IN1(n7053), .IN2(n6281), .IN3(\FIFO[50][3] ), .IN4(n6282), 
        .Q(n2934) );
  AO22X1 U4259 ( .IN1(n7042), .IN2(n6281), .IN3(\FIFO[50][4] ), .IN4(n6282), 
        .Q(n2935) );
  AO22X1 U4260 ( .IN1(n7031), .IN2(n6281), .IN3(\FIFO[50][5] ), .IN4(n6282), 
        .Q(n2936) );
  AO22X1 U4261 ( .IN1(n7020), .IN2(n6281), .IN3(\FIFO[50][6] ), .IN4(n6282), 
        .Q(n2937) );
  AO22X1 U4262 ( .IN1(n7009), .IN2(n6280), .IN3(\FIFO[50][7] ), .IN4(n6282), 
        .Q(n2938) );
  AO22X1 U4263 ( .IN1(n6998), .IN2(n6280), .IN3(\FIFO[50][8] ), .IN4(n6282), 
        .Q(n2939) );
  AO22X1 U4264 ( .IN1(n6987), .IN2(n6280), .IN3(\FIFO[50][9] ), .IN4(n6282), 
        .Q(n2940) );
  AO22X1 U4265 ( .IN1(n6976), .IN2(n6280), .IN3(\FIFO[50][10] ), .IN4(n6282), 
        .Q(n2941) );
  AO22X1 U4266 ( .IN1(n6965), .IN2(n6280), .IN3(\FIFO[50][11] ), .IN4(n6282), 
        .Q(n2942) );
  AO22X1 U4267 ( .IN1(n6954), .IN2(n6280), .IN3(\FIFO[50][12] ), .IN4(n6283), 
        .Q(n2943) );
  AO22X1 U4268 ( .IN1(n6943), .IN2(n6280), .IN3(\FIFO[50][13] ), .IN4(n6283), 
        .Q(n2944) );
  AO22X1 U4269 ( .IN1(n6932), .IN2(n6279), .IN3(\FIFO[50][14] ), .IN4(n6283), 
        .Q(n2945) );
  AO22X1 U4270 ( .IN1(n6921), .IN2(n6279), .IN3(\FIFO[50][15] ), .IN4(n6283), 
        .Q(n2946) );
  AO22X1 U4271 ( .IN1(n6910), .IN2(n6279), .IN3(\FIFO[50][16] ), .IN4(n6283), 
        .Q(n2947) );
  AO22X1 U4272 ( .IN1(n6899), .IN2(n6279), .IN3(\FIFO[50][17] ), .IN4(n6283), 
        .Q(n2948) );
  AO22X1 U4273 ( .IN1(n6888), .IN2(n6279), .IN3(\FIFO[50][18] ), .IN4(n6283), 
        .Q(n2949) );
  AO22X1 U4274 ( .IN1(n6877), .IN2(n6279), .IN3(\FIFO[50][19] ), .IN4(n6283), 
        .Q(n2950) );
  AO22X1 U4275 ( .IN1(n6866), .IN2(n6279), .IN3(\FIFO[50][20] ), .IN4(n6283), 
        .Q(n2951) );
  AO22X1 U4276 ( .IN1(n6855), .IN2(n6281), .IN3(\FIFO[50][21] ), .IN4(n6283), 
        .Q(n2952) );
  AO22X1 U4277 ( .IN1(n6844), .IN2(n6280), .IN3(\FIFO[50][22] ), .IN4(n6283), 
        .Q(n2953) );
  AO22X1 U4278 ( .IN1(n6833), .IN2(n6279), .IN3(\FIFO[50][23] ), .IN4(n6283), 
        .Q(n2954) );
  AO22X1 U4279 ( .IN1(n7091), .IN2(n6263), .IN3(\FIFO[47][0] ), .IN4(n6264), 
        .Q(n3027) );
  AO22X1 U4280 ( .IN1(n7074), .IN2(n6263), .IN3(\FIFO[47][1] ), .IN4(n6264), 
        .Q(n3028) );
  AO22X1 U4286 ( .IN1(n7063), .IN2(n6263), .IN3(\FIFO[47][2] ), .IN4(n6264), 
        .Q(n3029) );
  AO22X1 U4291 ( .IN1(n7052), .IN2(n6263), .IN3(\FIFO[47][3] ), .IN4(n6264), 
        .Q(n3030) );
  AO22X1 U4292 ( .IN1(n7041), .IN2(n6263), .IN3(\FIFO[47][4] ), .IN4(n6264), 
        .Q(n3031) );
  AO22X1 U4293 ( .IN1(n7030), .IN2(n6263), .IN3(\FIFO[47][5] ), .IN4(n6264), 
        .Q(n3032) );
  AO22X1 U4294 ( .IN1(n7019), .IN2(n6263), .IN3(\FIFO[47][6] ), .IN4(n6264), 
        .Q(n3033) );
  AO22X1 U4295 ( .IN1(n7008), .IN2(n6262), .IN3(\FIFO[47][7] ), .IN4(n6264), 
        .Q(n3034) );
  AO22X1 U4296 ( .IN1(n6997), .IN2(n6262), .IN3(\FIFO[47][8] ), .IN4(n6264), 
        .Q(n3035) );
  AO22X1 U4297 ( .IN1(n6986), .IN2(n6262), .IN3(\FIFO[47][9] ), .IN4(n6264), 
        .Q(n3036) );
  AO22X1 U4298 ( .IN1(n6975), .IN2(n6262), .IN3(\FIFO[47][10] ), .IN4(n6264), 
        .Q(n3037) );
  AO22X1 U4299 ( .IN1(n6964), .IN2(n6262), .IN3(\FIFO[47][11] ), .IN4(n6264), 
        .Q(n3038) );
  AO22X1 U4300 ( .IN1(n6953), .IN2(n6262), .IN3(\FIFO[47][12] ), .IN4(n6265), 
        .Q(n3039) );
  AO22X1 U4301 ( .IN1(n6942), .IN2(n6262), .IN3(\FIFO[47][13] ), .IN4(n6265), 
        .Q(n3040) );
  AO22X1 U4302 ( .IN1(n6931), .IN2(n6261), .IN3(\FIFO[47][14] ), .IN4(n6265), 
        .Q(n3041) );
  AO22X1 U4303 ( .IN1(n6920), .IN2(n6261), .IN3(\FIFO[47][15] ), .IN4(n6265), 
        .Q(n3042) );
  AO22X1 U4304 ( .IN1(n6909), .IN2(n6261), .IN3(\FIFO[47][16] ), .IN4(n6265), 
        .Q(n3043) );
  AO22X1 U4305 ( .IN1(n6898), .IN2(n6261), .IN3(\FIFO[47][17] ), .IN4(n6265), 
        .Q(n3044) );
  AO22X1 U4306 ( .IN1(n6887), .IN2(n6261), .IN3(\FIFO[47][18] ), .IN4(n6265), 
        .Q(n3045) );
  AO22X1 U4307 ( .IN1(n6876), .IN2(n6261), .IN3(\FIFO[47][19] ), .IN4(n6265), 
        .Q(n3046) );
  AO22X1 U4308 ( .IN1(n6865), .IN2(n6261), .IN3(\FIFO[47][20] ), .IN4(n6265), 
        .Q(n3047) );
  AO22X1 U4309 ( .IN1(n6854), .IN2(n6263), .IN3(\FIFO[47][21] ), .IN4(n6265), 
        .Q(n3048) );
  AO22X1 U4310 ( .IN1(n6843), .IN2(n6262), .IN3(\FIFO[47][22] ), .IN4(n6265), 
        .Q(n3049) );
  AO22X1 U4311 ( .IN1(n6832), .IN2(n6261), .IN3(\FIFO[47][23] ), .IN4(n6265), 
        .Q(n3050) );
  AO22X1 U4312 ( .IN1(n7091), .IN2(n6257), .IN3(\FIFO[46][0] ), .IN4(n6258), 
        .Q(n3059) );
  AO22X1 U4313 ( .IN1(n7074), .IN2(n6257), .IN3(\FIFO[46][1] ), .IN4(n6258), 
        .Q(n3060) );
  AO22X1 U4314 ( .IN1(n7063), .IN2(n6257), .IN3(\FIFO[46][2] ), .IN4(n6258), 
        .Q(n3061) );
  AO22X1 U4323 ( .IN1(n7052), .IN2(n6257), .IN3(\FIFO[46][3] ), .IN4(n6258), 
        .Q(n3062) );
  AO22X1 U4324 ( .IN1(n7041), .IN2(n6257), .IN3(\FIFO[46][4] ), .IN4(n6258), 
        .Q(n3063) );
  AO22X1 U4334 ( .IN1(n7030), .IN2(n6257), .IN3(\FIFO[46][5] ), .IN4(n6258), 
        .Q(n3064) );
  AO22X1 U4345 ( .IN1(n7019), .IN2(n6257), .IN3(\FIFO[46][6] ), .IN4(n6258), 
        .Q(n3065) );
  AO22X1 U4357 ( .IN1(n7008), .IN2(n6256), .IN3(\FIFO[46][7] ), .IN4(n6258), 
        .Q(n3066) );
  AO22X1 U4358 ( .IN1(n6997), .IN2(n6256), .IN3(\FIFO[46][8] ), .IN4(n6258), 
        .Q(n3067) );
  AO22X1 U4369 ( .IN1(n6986), .IN2(n6256), .IN3(\FIFO[46][9] ), .IN4(n6258), 
        .Q(n3068) );
  AO22X1 U4380 ( .IN1(n6975), .IN2(n6256), .IN3(\FIFO[46][10] ), .IN4(n6258), 
        .Q(n3069) );
  AO22X1 U4393 ( .IN1(n6964), .IN2(n6256), .IN3(\FIFO[46][11] ), .IN4(n6258), 
        .Q(n3070) );
  AO22X1 U4394 ( .IN1(n6953), .IN2(n6256), .IN3(\FIFO[46][12] ), .IN4(n6259), 
        .Q(n3071) );
  AO22X1 U4395 ( .IN1(n6942), .IN2(n6256), .IN3(\FIFO[46][13] ), .IN4(n6259), 
        .Q(n3072) );
  AO22X1 U4396 ( .IN1(n6931), .IN2(n6255), .IN3(\FIFO[46][14] ), .IN4(n6259), 
        .Q(n3073) );
  AO22X1 U4397 ( .IN1(n6920), .IN2(n6255), .IN3(\FIFO[46][15] ), .IN4(n6259), 
        .Q(n3074) );
  AO22X1 U4398 ( .IN1(n6909), .IN2(n6255), .IN3(\FIFO[46][16] ), .IN4(n6259), 
        .Q(n3075) );
  AO22X1 U4399 ( .IN1(n6898), .IN2(n6255), .IN3(\FIFO[46][17] ), .IN4(n6259), 
        .Q(n3076) );
  AO22X1 U4400 ( .IN1(n6887), .IN2(n6255), .IN3(\FIFO[46][18] ), .IN4(n6259), 
        .Q(n3077) );
  AO22X1 U4401 ( .IN1(n6876), .IN2(n6255), .IN3(\FIFO[46][19] ), .IN4(n6259), 
        .Q(n3078) );
  AO22X1 U4402 ( .IN1(n6865), .IN2(n6255), .IN3(\FIFO[46][20] ), .IN4(n6259), 
        .Q(n3079) );
  AO22X1 U4403 ( .IN1(n6854), .IN2(n6257), .IN3(\FIFO[46][21] ), .IN4(n6259), 
        .Q(n3080) );
  AO22X1 U4404 ( .IN1(n6843), .IN2(n6256), .IN3(\FIFO[46][22] ), .IN4(n6259), 
        .Q(n3081) );
  AO22X1 U4405 ( .IN1(n6832), .IN2(n6255), .IN3(\FIFO[46][23] ), .IN4(n6259), 
        .Q(n3082) );
  AO22X1 U4406 ( .IN1(n7091), .IN2(n6239), .IN3(\FIFO[43][0] ), .IN4(n6240), 
        .Q(n3155) );
  AO22X1 U4407 ( .IN1(n7063), .IN2(n6237), .IN3(\FIFO[43][2] ), .IN4(n6240), 
        .Q(n3157) );
  AO22X1 U4408 ( .IN1(n7052), .IN2(n6239), .IN3(\FIFO[43][3] ), .IN4(n6240), 
        .Q(n3158) );
  AO22X1 U4409 ( .IN1(n7041), .IN2(n6238), .IN3(\FIFO[43][4] ), .IN4(n6240), 
        .Q(n3159) );
  AO22X1 U4410 ( .IN1(n7030), .IN2(n6237), .IN3(\FIFO[43][5] ), .IN4(n6240), 
        .Q(n3160) );
  AO22X1 U4411 ( .IN1(n7019), .IN2(n6239), .IN3(\FIFO[43][6] ), .IN4(n6240), 
        .Q(n3161) );
  AO22X1 U4412 ( .IN1(n7008), .IN2(n6239), .IN3(\FIFO[43][7] ), .IN4(n6240), 
        .Q(n3162) );
  AO22X1 U4413 ( .IN1(n6997), .IN2(n6239), .IN3(\FIFO[43][8] ), .IN4(n6240), 
        .Q(n3163) );
  AO22X1 U4414 ( .IN1(n6986), .IN2(n6239), .IN3(\FIFO[43][9] ), .IN4(n6240), 
        .Q(n3164) );
  AO22X1 U4415 ( .IN1(n6975), .IN2(n6239), .IN3(\FIFO[43][10] ), .IN4(n6240), 
        .Q(n3165) );
  AO22X1 U4416 ( .IN1(n6964), .IN2(n6239), .IN3(\FIFO[43][11] ), .IN4(n6240), 
        .Q(n3166) );
  AO22X1 U4423 ( .IN1(n6953), .IN2(n6239), .IN3(\FIFO[43][12] ), .IN4(n6241), 
        .Q(n3167) );
  AO22X1 U4427 ( .IN1(n6942), .IN2(n6239), .IN3(\FIFO[43][13] ), .IN4(n6241), 
        .Q(n3168) );
  AO22X1 U4428 ( .IN1(n6931), .IN2(n6238), .IN3(\FIFO[43][14] ), .IN4(n6241), 
        .Q(n3169) );
  AO22X1 U4429 ( .IN1(n6920), .IN2(n6238), .IN3(\FIFO[43][15] ), .IN4(n6241), 
        .Q(n3170) );
  AO22X1 U4430 ( .IN1(n6909), .IN2(n6238), .IN3(\FIFO[43][16] ), .IN4(n6241), 
        .Q(n3171) );
  AO22X1 U4431 ( .IN1(n6898), .IN2(n6238), .IN3(\FIFO[43][17] ), .IN4(n6241), 
        .Q(n3172) );
  AO22X1 U4432 ( .IN1(n6887), .IN2(n6238), .IN3(\FIFO[43][18] ), .IN4(n6241), 
        .Q(n3173) );
  AO22X1 U4433 ( .IN1(n6876), .IN2(n6238), .IN3(\FIFO[43][19] ), .IN4(n6241), 
        .Q(n3174) );
  AO22X1 U4434 ( .IN1(n6865), .IN2(n6238), .IN3(\FIFO[43][20] ), .IN4(n6241), 
        .Q(n3175) );
  AO22X1 U4435 ( .IN1(n6854), .IN2(n6237), .IN3(\FIFO[43][21] ), .IN4(n6241), 
        .Q(n3176) );
  AO22X1 U4436 ( .IN1(n6832), .IN2(n6237), .IN3(\FIFO[43][23] ), .IN4(n6241), 
        .Q(n3178) );
  AO22X1 U4437 ( .IN1(n7091), .IN2(n6233), .IN3(\FIFO[42][0] ), .IN4(n6234), 
        .Q(n3187) );
  AO22X1 U4438 ( .IN1(n7074), .IN2(n6233), .IN3(\FIFO[42][1] ), .IN4(n6234), 
        .Q(n3188) );
  AO22X1 U4439 ( .IN1(n7063), .IN2(n6233), .IN3(\FIFO[42][2] ), .IN4(n6234), 
        .Q(n3189) );
  AO22X1 U4440 ( .IN1(n7052), .IN2(n6233), .IN3(\FIFO[42][3] ), .IN4(n6234), 
        .Q(n3190) );
  AO22X1 U4441 ( .IN1(n7030), .IN2(n6233), .IN3(\FIFO[42][5] ), .IN4(n6234), 
        .Q(n3192) );
  AO22X1 U4442 ( .IN1(n7019), .IN2(n6233), .IN3(\FIFO[42][6] ), .IN4(n6234), 
        .Q(n3193) );
  AO22X1 U4443 ( .IN1(n7008), .IN2(n6232), .IN3(\FIFO[42][7] ), .IN4(n6234), 
        .Q(n3194) );
  AO22X1 U4444 ( .IN1(n6997), .IN2(n6232), .IN3(\FIFO[42][8] ), .IN4(n6234), 
        .Q(n3195) );
  AO22X1 U4445 ( .IN1(n6986), .IN2(n6232), .IN3(\FIFO[42][9] ), .IN4(n6234), 
        .Q(n3196) );
  AO22X1 U4446 ( .IN1(n6975), .IN2(n6232), .IN3(\FIFO[42][10] ), .IN4(n6234), 
        .Q(n3197) );
  AO22X1 U4447 ( .IN1(n6964), .IN2(n6232), .IN3(\FIFO[42][11] ), .IN4(n6234), 
        .Q(n3198) );
  AO22X1 U4448 ( .IN1(n6953), .IN2(n6232), .IN3(\FIFO[42][12] ), .IN4(n6235), 
        .Q(n3199) );
  AO22X1 U4449 ( .IN1(n6942), .IN2(n6232), .IN3(\FIFO[42][13] ), .IN4(n6235), 
        .Q(n3200) );
  AO22X1 U4450 ( .IN1(n6931), .IN2(n6231), .IN3(\FIFO[42][14] ), .IN4(n6235), 
        .Q(n3201) );
  AO22X1 U4458 ( .IN1(n6920), .IN2(n6231), .IN3(\FIFO[42][15] ), .IN4(n6235), 
        .Q(n3202) );
  AO22X1 U4467 ( .IN1(n6909), .IN2(n6231), .IN3(\FIFO[42][16] ), .IN4(n6235), 
        .Q(n3203) );
  AO22X1 U4483 ( .IN1(n6898), .IN2(n6231), .IN3(\FIFO[42][17] ), .IN4(n6235), 
        .Q(n3204) );
  AO22X1 U4496 ( .IN1(n6887), .IN2(n6231), .IN3(\FIFO[42][18] ), .IN4(n6235), 
        .Q(n3205) );
  AO22X1 U4498 ( .IN1(n6876), .IN2(n6231), .IN3(\FIFO[42][19] ), .IN4(n6235), 
        .Q(n3206) );
  AO22X1 U4500 ( .IN1(n6865), .IN2(n6231), .IN3(\FIFO[42][20] ), .IN4(n6235), 
        .Q(n3207) );
  AO22X1 U4502 ( .IN1(n6854), .IN2(n6233), .IN3(\FIFO[42][21] ), .IN4(n6235), 
        .Q(n3208) );
  AO22X1 U4504 ( .IN1(n6843), .IN2(n6232), .IN3(\FIFO[42][22] ), .IN4(n6235), 
        .Q(n3209) );
  AO22X1 U4506 ( .IN1(n6832), .IN2(n6231), .IN3(\FIFO[42][23] ), .IN4(n6235), 
        .Q(n3210) );
  AO22X1 U4508 ( .IN1(n7091), .IN2(n6215), .IN3(\FIFO[39][0] ), .IN4(n6216), 
        .Q(n3283) );
  AO22X1 U4510 ( .IN1(n7074), .IN2(n6215), .IN3(\FIFO[39][1] ), .IN4(n6216), 
        .Q(n3284) );
  AO22X1 U4512 ( .IN1(n7063), .IN2(n6215), .IN3(\FIFO[39][2] ), .IN4(n6216), 
        .Q(n3285) );
  AO22X1 U4514 ( .IN1(n7052), .IN2(n6215), .IN3(\FIFO[39][3] ), .IN4(n6216), 
        .Q(n3286) );
  AO22X1 U4516 ( .IN1(n7041), .IN2(n6215), .IN3(\FIFO[39][4] ), .IN4(n6216), 
        .Q(n3287) );
  AO22X1 U4517 ( .IN1(n7030), .IN2(n6215), .IN3(\FIFO[39][5] ), .IN4(n6216), 
        .Q(n3288) );
  AO22X1 U4518 ( .IN1(n7019), .IN2(n6215), .IN3(\FIFO[39][6] ), .IN4(n6216), 
        .Q(n3289) );
  AO22X1 U4520 ( .IN1(n7008), .IN2(n6214), .IN3(\FIFO[39][7] ), .IN4(n6216), 
        .Q(n3290) );
  AO22X1 U4522 ( .IN1(n6997), .IN2(n6214), .IN3(\FIFO[39][8] ), .IN4(n6216), 
        .Q(n3291) );
  AO22X1 U4524 ( .IN1(n6986), .IN2(n6214), .IN3(\FIFO[39][9] ), .IN4(n6216), 
        .Q(n3292) );
  AO22X1 U4526 ( .IN1(n6975), .IN2(n6214), .IN3(\FIFO[39][10] ), .IN4(n6216), 
        .Q(n3293) );
  AO22X1 U4528 ( .IN1(n6964), .IN2(n6214), .IN3(\FIFO[39][11] ), .IN4(n6216), 
        .Q(n3294) );
  AO22X1 U4530 ( .IN1(n6953), .IN2(n6214), .IN3(\FIFO[39][12] ), .IN4(n6217), 
        .Q(n3295) );
  AO22X1 U4532 ( .IN1(n6942), .IN2(n6214), .IN3(\FIFO[39][13] ), .IN4(n6217), 
        .Q(n3296) );
  AO22X1 U4534 ( .IN1(n6920), .IN2(n6214), .IN3(\FIFO[39][15] ), .IN4(n6217), 
        .Q(n3298) );
  AO22X1 U4536 ( .IN1(n6909), .IN2(n6213), .IN3(\FIFO[39][16] ), .IN4(n6217), 
        .Q(n3299) );
  AO22X1 U4538 ( .IN1(n6898), .IN2(n6215), .IN3(\FIFO[39][17] ), .IN4(n6217), 
        .Q(n3300) );
  AO22X1 U4540 ( .IN1(n6887), .IN2(n6214), .IN3(\FIFO[39][18] ), .IN4(n6217), 
        .Q(n3301) );
  AO22X1 U4541 ( .IN1(n6876), .IN2(n6213), .IN3(\FIFO[39][19] ), .IN4(n6217), 
        .Q(n3302) );
  AO22X1 U4542 ( .IN1(n6865), .IN2(n6215), .IN3(\FIFO[39][20] ), .IN4(n6217), 
        .Q(n3303) );
  AO22X1 U4544 ( .IN1(n6854), .IN2(n6213), .IN3(\FIFO[39][21] ), .IN4(n6217), 
        .Q(n3304) );
  AO22X1 U4546 ( .IN1(n6843), .IN2(n6213), .IN3(\FIFO[39][22] ), .IN4(n6217), 
        .Q(n3305) );
  AO22X1 U4548 ( .IN1(n7091), .IN2(n6209), .IN3(\FIFO[38][0] ), .IN4(n6210), 
        .Q(n3315) );
  AO22X1 U4550 ( .IN1(n7074), .IN2(n6208), .IN3(\FIFO[38][1] ), .IN4(n6210), 
        .Q(n3316) );
  AO22X1 U4552 ( .IN1(n7063), .IN2(n6207), .IN3(\FIFO[38][2] ), .IN4(n6210), 
        .Q(n3317) );
  AO22X1 U4554 ( .IN1(n7052), .IN2(n6209), .IN3(\FIFO[38][3] ), .IN4(n6210), 
        .Q(n3318) );
  AO22X1 U4556 ( .IN1(n7041), .IN2(n6208), .IN3(\FIFO[38][4] ), .IN4(n6210), 
        .Q(n3319) );
  AO22X1 U4560 ( .IN1(n7030), .IN2(n6207), .IN3(\FIFO[38][5] ), .IN4(n6210), 
        .Q(n3320) );
  AO22X1 U4561 ( .IN1(n7019), .IN2(n6209), .IN3(\FIFO[38][6] ), .IN4(n6210), 
        .Q(n3321) );
  AO22X1 U4562 ( .IN1(n7008), .IN2(n6209), .IN3(\FIFO[38][7] ), .IN4(n6210), 
        .Q(n3322) );
  AO22X1 U4563 ( .IN1(n6997), .IN2(n6209), .IN3(\FIFO[38][8] ), .IN4(n6210), 
        .Q(n3323) );
  AO22X1 U4564 ( .IN1(n6986), .IN2(n6209), .IN3(\FIFO[38][9] ), .IN4(n6210), 
        .Q(n3324) );
  AO22X1 U4593 ( .IN1(n6975), .IN2(n6209), .IN3(\FIFO[38][10] ), .IN4(n6210), 
        .Q(n3325) );
  AO22X1 U4596 ( .IN1(n6964), .IN2(n6209), .IN3(\FIFO[38][11] ), .IN4(n6210), 
        .Q(n3326) );
  AO22X1 U4597 ( .IN1(n6953), .IN2(n6209), .IN3(\FIFO[38][12] ), .IN4(n6211), 
        .Q(n3327) );
  AO22X1 U4598 ( .IN1(n6942), .IN2(n6209), .IN3(\FIFO[38][13] ), .IN4(n6211), 
        .Q(n3328) );
  AO22X1 U4599 ( .IN1(n6931), .IN2(n6208), .IN3(\FIFO[38][14] ), .IN4(n6211), 
        .Q(n3329) );
  AO22X1 U4600 ( .IN1(n6920), .IN2(n6208), .IN3(\FIFO[38][15] ), .IN4(n6211), 
        .Q(n3330) );
  AO22X1 U4601 ( .IN1(n6898), .IN2(n6208), .IN3(\FIFO[38][17] ), .IN4(n6211), 
        .Q(n3332) );
  AO22X1 U4602 ( .IN1(n6887), .IN2(n6208), .IN3(\FIFO[38][18] ), .IN4(n6211), 
        .Q(n3333) );
  AO22X1 U4603 ( .IN1(n6876), .IN2(n6208), .IN3(\FIFO[38][19] ), .IN4(n6211), 
        .Q(n3334) );
  AO22X1 U4604 ( .IN1(n6865), .IN2(n6208), .IN3(\FIFO[38][20] ), .IN4(n6211), 
        .Q(n3335) );
  AO22X1 U4605 ( .IN1(n6854), .IN2(n6207), .IN3(\FIFO[38][21] ), .IN4(n6211), 
        .Q(n3336) );
  AO22X1 U4606 ( .IN1(n6843), .IN2(n6207), .IN3(\FIFO[38][22] ), .IN4(n6211), 
        .Q(n3337) );
  AO22X1 U4607 ( .IN1(n6832), .IN2(n6207), .IN3(\FIFO[38][23] ), .IN4(n6211), 
        .Q(n3338) );
  AO22X1 U4608 ( .IN1(n7090), .IN2(n6191), .IN3(\FIFO[35][0] ), .IN4(n6192), 
        .Q(n3411) );
  AO22X1 U4609 ( .IN1(n7073), .IN2(n6191), .IN3(\FIFO[35][1] ), .IN4(n6192), 
        .Q(n3412) );
  AO22X1 U4610 ( .IN1(n7062), .IN2(n6191), .IN3(\FIFO[35][2] ), .IN4(n6192), 
        .Q(n3413) );
  AO22X1 U4611 ( .IN1(n7051), .IN2(n6191), .IN3(\FIFO[35][3] ), .IN4(n6192), 
        .Q(n3414) );
  AO22X1 U4612 ( .IN1(n7040), .IN2(n6191), .IN3(\FIFO[35][4] ), .IN4(n6192), 
        .Q(n3415) );
  AO22X1 U4613 ( .IN1(n7029), .IN2(n6191), .IN3(\FIFO[35][5] ), .IN4(n6192), 
        .Q(n3416) );
  AO22X1 U4614 ( .IN1(n7018), .IN2(n6191), .IN3(\FIFO[35][6] ), .IN4(n6192), 
        .Q(n3417) );
  AO22X1 U4615 ( .IN1(n7007), .IN2(n6190), .IN3(\FIFO[35][7] ), .IN4(n6192), 
        .Q(n3418) );
  AO22X1 U4616 ( .IN1(n6996), .IN2(n6190), .IN3(\FIFO[35][8] ), .IN4(n6192), 
        .Q(n3419) );
  AO22X1 U4617 ( .IN1(n6985), .IN2(n6190), .IN3(\FIFO[35][9] ), .IN4(n6192), 
        .Q(n3420) );
  AO22X1 U4618 ( .IN1(n6974), .IN2(n6190), .IN3(\FIFO[35][10] ), .IN4(n6192), 
        .Q(n3421) );
  AO22X1 U4619 ( .IN1(n6963), .IN2(n6190), .IN3(\FIFO[35][11] ), .IN4(n6192), 
        .Q(n3422) );
  AO22X1 U4620 ( .IN1(n6952), .IN2(n6190), .IN3(\FIFO[35][12] ), .IN4(n6193), 
        .Q(n3423) );
  AO22X1 U4621 ( .IN1(n6941), .IN2(n6190), .IN3(\FIFO[35][13] ), .IN4(n6193), 
        .Q(n3424) );
  AO22X1 U4622 ( .IN1(n6919), .IN2(n6189), .IN3(\FIFO[35][15] ), .IN4(n6193), 
        .Q(n3426) );
  AO22X1 U4623 ( .IN1(n6908), .IN2(n6189), .IN3(\FIFO[35][16] ), .IN4(n6193), 
        .Q(n3427) );
  AO22X1 U4624 ( .IN1(n6897), .IN2(n6189), .IN3(\FIFO[35][17] ), .IN4(n6193), 
        .Q(n3428) );
  AO22X1 U4625 ( .IN1(n6886), .IN2(n6189), .IN3(\FIFO[35][18] ), .IN4(n6193), 
        .Q(n3429) );
  AO22X1 U4626 ( .IN1(n6875), .IN2(n6189), .IN3(\FIFO[35][19] ), .IN4(n6193), 
        .Q(n3430) );
  AO22X1 U4627 ( .IN1(n6864), .IN2(n6189), .IN3(\FIFO[35][20] ), .IN4(n6193), 
        .Q(n3431) );
  AO22X1 U4628 ( .IN1(n6853), .IN2(n6191), .IN3(\FIFO[35][21] ), .IN4(n6193), 
        .Q(n3432) );
  AO22X1 U4629 ( .IN1(n6842), .IN2(n6190), .IN3(\FIFO[35][22] ), .IN4(n6193), 
        .Q(n3433) );
  AO22X1 U4630 ( .IN1(n6831), .IN2(n6189), .IN3(\FIFO[35][23] ), .IN4(n6193), 
        .Q(n3434) );
  AO22X1 U4631 ( .IN1(n7090), .IN2(n6185), .IN3(\FIFO[34][0] ), .IN4(n6186), 
        .Q(n3443) );
  AO22X1 U4632 ( .IN1(n7073), .IN2(n6185), .IN3(\FIFO[34][1] ), .IN4(n6186), 
        .Q(n3444) );
  AO22X1 U4633 ( .IN1(n7062), .IN2(n6185), .IN3(\FIFO[34][2] ), .IN4(n6186), 
        .Q(n3445) );
  AO22X1 U4634 ( .IN1(n7051), .IN2(n6185), .IN3(\FIFO[34][3] ), .IN4(n6186), 
        .Q(n3446) );
  AO22X1 U4635 ( .IN1(n7040), .IN2(n6185), .IN3(\FIFO[34][4] ), .IN4(n6186), 
        .Q(n3447) );
  AO22X1 U4636 ( .IN1(n7029), .IN2(n6185), .IN3(\FIFO[34][5] ), .IN4(n6186), 
        .Q(n3448) );
  AO22X1 U4637 ( .IN1(n7018), .IN2(n6185), .IN3(\FIFO[34][6] ), .IN4(n6186), 
        .Q(n3449) );
  AO22X1 U4638 ( .IN1(n7007), .IN2(n6184), .IN3(\FIFO[34][7] ), .IN4(n6186), 
        .Q(n3450) );
  AO22X1 U4639 ( .IN1(n6996), .IN2(n6184), .IN3(\FIFO[34][8] ), .IN4(n6186), 
        .Q(n3451) );
  AO22X1 U4640 ( .IN1(n6985), .IN2(n6184), .IN3(\FIFO[34][9] ), .IN4(n6186), 
        .Q(n3452) );
  AO22X1 U4641 ( .IN1(n6974), .IN2(n6184), .IN3(\FIFO[34][10] ), .IN4(n6186), 
        .Q(n3453) );
  AO22X1 U4642 ( .IN1(n6952), .IN2(n6184), .IN3(\FIFO[34][12] ), .IN4(n6187), 
        .Q(n3455) );
  AO22X1 U4643 ( .IN1(n6941), .IN2(n6184), .IN3(\FIFO[34][13] ), .IN4(n6187), 
        .Q(n3456) );
  AO22X1 U4644 ( .IN1(n6930), .IN2(n6185), .IN3(\FIFO[34][14] ), .IN4(n6187), 
        .Q(n3457) );
  AO22X1 U4645 ( .IN1(n6919), .IN2(n6184), .IN3(\FIFO[34][15] ), .IN4(n6187), 
        .Q(n3458) );
  AO22X1 U4646 ( .IN1(n6908), .IN2(n6183), .IN3(\FIFO[34][16] ), .IN4(n6187), 
        .Q(n3459) );
  AO22X1 U4647 ( .IN1(n6886), .IN2(n6184), .IN3(\FIFO[34][18] ), .IN4(n6187), 
        .Q(n3461) );
  AO22X1 U4648 ( .IN1(n6875), .IN2(n6183), .IN3(\FIFO[34][19] ), .IN4(n6187), 
        .Q(n3462) );
  AO22X1 U4649 ( .IN1(n6864), .IN2(n6185), .IN3(\FIFO[34][20] ), .IN4(n6187), 
        .Q(n3463) );
  AO22X1 U4650 ( .IN1(n6853), .IN2(n6183), .IN3(\FIFO[34][21] ), .IN4(n6187), 
        .Q(n3464) );
  AO22X1 U4651 ( .IN1(n6842), .IN2(n6183), .IN3(\FIFO[34][22] ), .IN4(n6187), 
        .Q(n3465) );
  AO22X1 U4652 ( .IN1(n6831), .IN2(n6183), .IN3(\FIFO[34][23] ), .IN4(n6187), 
        .Q(n3466) );
  AO22X1 U4653 ( .IN1(n7073), .IN2(n6166), .IN3(\FIFO[31][1] ), .IN4(n6168), 
        .Q(n3540) );
  AO22X1 U4654 ( .IN1(n7062), .IN2(n6165), .IN3(\FIFO[31][2] ), .IN4(n6168), 
        .Q(n3541) );
  AO22X1 U4655 ( .IN1(n7051), .IN2(n6167), .IN3(\FIFO[31][3] ), .IN4(n6168), 
        .Q(n3542) );
  AO22X1 U4656 ( .IN1(n7040), .IN2(n6166), .IN3(\FIFO[31][4] ), .IN4(n6168), 
        .Q(n3543) );
  AO22X1 U4657 ( .IN1(n7029), .IN2(n6165), .IN3(\FIFO[31][5] ), .IN4(n6168), 
        .Q(n3544) );
  AO22X1 U4658 ( .IN1(n7018), .IN2(n6167), .IN3(\FIFO[31][6] ), .IN4(n6168), 
        .Q(n3545) );
  AO22X1 U4659 ( .IN1(n7007), .IN2(n6167), .IN3(\FIFO[31][7] ), .IN4(n6168), 
        .Q(n3546) );
  AO22X1 U4660 ( .IN1(n6996), .IN2(n6167), .IN3(\FIFO[31][8] ), .IN4(n6168), 
        .Q(n3547) );
  AO22X1 U4661 ( .IN1(n6985), .IN2(n6167), .IN3(\FIFO[31][9] ), .IN4(n6168), 
        .Q(n3548) );
  AO22X1 U4662 ( .IN1(n6974), .IN2(n6167), .IN3(\FIFO[31][10] ), .IN4(n6168), 
        .Q(n3549) );
  AO22X1 U4663 ( .IN1(n6963), .IN2(n6167), .IN3(\FIFO[31][11] ), .IN4(n6168), 
        .Q(n3550) );
  AO22X1 U4664 ( .IN1(n6952), .IN2(n6167), .IN3(\FIFO[31][12] ), .IN4(n6169), 
        .Q(n3551) );
  AO22X1 U4665 ( .IN1(n6941), .IN2(n6167), .IN3(\FIFO[31][13] ), .IN4(n6169), 
        .Q(n3552) );
  AO22X1 U4666 ( .IN1(n6930), .IN2(n6166), .IN3(\FIFO[31][14] ), .IN4(n6169), 
        .Q(n3553) );
  AO22X1 U4667 ( .IN1(n6919), .IN2(n6166), .IN3(\FIFO[31][15] ), .IN4(n6169), 
        .Q(n3554) );
  AO22X1 U4668 ( .IN1(n6908), .IN2(n6166), .IN3(\FIFO[31][16] ), .IN4(n6169), 
        .Q(n3555) );
  AO22X1 U4669 ( .IN1(n6897), .IN2(n6166), .IN3(\FIFO[31][17] ), .IN4(n6169), 
        .Q(n3556) );
  AO22X1 U4670 ( .IN1(n6886), .IN2(n6166), .IN3(\FIFO[31][18] ), .IN4(n6169), 
        .Q(n3557) );
  AO22X1 U4671 ( .IN1(n6864), .IN2(n6166), .IN3(\FIFO[31][20] ), .IN4(n6169), 
        .Q(n3559) );
  AO22X1 U4672 ( .IN1(n6853), .IN2(n6165), .IN3(\FIFO[31][21] ), .IN4(n6169), 
        .Q(n3560) );
  AO22X1 U4673 ( .IN1(n6842), .IN2(n6165), .IN3(\FIFO[31][22] ), .IN4(n6169), 
        .Q(n3561) );
  AO22X1 U4674 ( .IN1(n6831), .IN2(n6165), .IN3(\FIFO[31][23] ), .IN4(n6169), 
        .Q(n3562) );
  AO22X1 U4675 ( .IN1(n7090), .IN2(n6161), .IN3(\FIFO[30][0] ), .IN4(n6162), 
        .Q(n3571) );
  AO22X1 U4676 ( .IN1(n7062), .IN2(n6161), .IN3(\FIFO[30][2] ), .IN4(n6162), 
        .Q(n3573) );
  AO22X1 U4677 ( .IN1(n7051), .IN2(n6161), .IN3(\FIFO[30][3] ), .IN4(n6162), 
        .Q(n3574) );
  AO22X1 U4678 ( .IN1(n7040), .IN2(n6161), .IN3(\FIFO[30][4] ), .IN4(n6162), 
        .Q(n3575) );
  AO22X1 U4679 ( .IN1(n7029), .IN2(n6161), .IN3(\FIFO[30][5] ), .IN4(n6162), 
        .Q(n3576) );
  AO22X1 U4680 ( .IN1(n7018), .IN2(n6161), .IN3(\FIFO[30][6] ), .IN4(n6162), 
        .Q(n3577) );
  AO22X1 U4681 ( .IN1(n7007), .IN2(n6160), .IN3(\FIFO[30][7] ), .IN4(n6162), 
        .Q(n3578) );
  AO22X1 U4682 ( .IN1(n6996), .IN2(n6160), .IN3(\FIFO[30][8] ), .IN4(n6162), 
        .Q(n3579) );
  AO22X1 U4683 ( .IN1(n6985), .IN2(n6160), .IN3(\FIFO[30][9] ), .IN4(n6162), 
        .Q(n3580) );
  AO22X1 U4684 ( .IN1(n6974), .IN2(n6160), .IN3(\FIFO[30][10] ), .IN4(n6162), 
        .Q(n3581) );
  AO22X1 U4685 ( .IN1(n6963), .IN2(n6160), .IN3(\FIFO[30][11] ), .IN4(n6162), 
        .Q(n3582) );
  AO22X1 U4686 ( .IN1(n6952), .IN2(n6160), .IN3(\FIFO[30][12] ), .IN4(n6163), 
        .Q(n3583) );
  AO22X1 U4687 ( .IN1(n6941), .IN2(n6160), .IN3(\FIFO[30][13] ), .IN4(n6163), 
        .Q(n3584) );
  AO22X1 U4688 ( .IN1(n6930), .IN2(n6159), .IN3(\FIFO[30][14] ), .IN4(n6163), 
        .Q(n3585) );
  AO22X1 U4689 ( .IN1(n6919), .IN2(n6159), .IN3(\FIFO[30][15] ), .IN4(n6163), 
        .Q(n3586) );
  AO22X1 U4690 ( .IN1(n6908), .IN2(n6159), .IN3(\FIFO[30][16] ), .IN4(n6163), 
        .Q(n3587) );
  AO22X1 U4691 ( .IN1(n6897), .IN2(n6159), .IN3(\FIFO[30][17] ), .IN4(n6163), 
        .Q(n3588) );
  AO22X1 U4692 ( .IN1(n6886), .IN2(n6159), .IN3(\FIFO[30][18] ), .IN4(n6163), 
        .Q(n3589) );
  AO22X1 U4693 ( .IN1(n6875), .IN2(n6159), .IN3(\FIFO[30][19] ), .IN4(n6163), 
        .Q(n3590) );
  AO22X1 U4694 ( .IN1(n6864), .IN2(n6159), .IN3(\FIFO[30][20] ), .IN4(n6163), 
        .Q(n3591) );
  AO22X1 U4695 ( .IN1(n6853), .IN2(n6161), .IN3(\FIFO[30][21] ), .IN4(n6163), 
        .Q(n3592) );
  AO22X1 U4696 ( .IN1(n6842), .IN2(n6160), .IN3(\FIFO[30][22] ), .IN4(n6163), 
        .Q(n3593) );
  AO22X1 U4697 ( .IN1(n6831), .IN2(n6159), .IN3(\FIFO[30][23] ), .IN4(n6163), 
        .Q(n3594) );
  AO22X1 U4698 ( .IN1(n7090), .IN2(n6143), .IN3(\FIFO[27][0] ), .IN4(n6144), 
        .Q(n3667) );
  AO22X1 U4699 ( .IN1(n7073), .IN2(n6143), .IN3(\FIFO[27][1] ), .IN4(n6144), 
        .Q(n3668) );
  AO22X1 U4700 ( .IN1(n7062), .IN2(n6143), .IN3(\FIFO[27][2] ), .IN4(n6144), 
        .Q(n3669) );
  AO22X1 U4701 ( .IN1(n7051), .IN2(n6143), .IN3(\FIFO[27][3] ), .IN4(n6144), 
        .Q(n3670) );
  AO22X1 U4702 ( .IN1(n7029), .IN2(n6143), .IN3(\FIFO[27][5] ), .IN4(n6144), 
        .Q(n3672) );
  AO22X1 U4703 ( .IN1(n7018), .IN2(n6143), .IN3(\FIFO[27][6] ), .IN4(n6144), 
        .Q(n3673) );
  AO22X1 U4704 ( .IN1(n7007), .IN2(n6142), .IN3(\FIFO[27][7] ), .IN4(n6144), 
        .Q(n3674) );
  AO22X1 U4705 ( .IN1(n6996), .IN2(n6142), .IN3(\FIFO[27][8] ), .IN4(n6144), 
        .Q(n3675) );
  AO22X1 U4706 ( .IN1(n6985), .IN2(n6142), .IN3(\FIFO[27][9] ), .IN4(n6144), 
        .Q(n3676) );
  AO22X1 U4707 ( .IN1(n6974), .IN2(n6142), .IN3(\FIFO[27][10] ), .IN4(n6144), 
        .Q(n3677) );
  AO22X1 U4708 ( .IN1(n6963), .IN2(n6142), .IN3(\FIFO[27][11] ), .IN4(n6144), 
        .Q(n3678) );
  AO22X1 U4709 ( .IN1(n6952), .IN2(n6142), .IN3(\FIFO[27][12] ), .IN4(n6145), 
        .Q(n3679) );
  AO22X1 U4710 ( .IN1(n6941), .IN2(n6142), .IN3(\FIFO[27][13] ), .IN4(n6145), 
        .Q(n3680) );
  AO22X1 U4711 ( .IN1(n6930), .IN2(n6143), .IN3(\FIFO[27][14] ), .IN4(n6145), 
        .Q(n3681) );
  AO22X1 U4712 ( .IN1(n6919), .IN2(n6142), .IN3(\FIFO[27][15] ), .IN4(n6145), 
        .Q(n3682) );
  AO22X1 U4713 ( .IN1(n6908), .IN2(n6141), .IN3(\FIFO[27][16] ), .IN4(n6145), 
        .Q(n3683) );
  AO22X1 U4714 ( .IN1(n6897), .IN2(n6143), .IN3(\FIFO[27][17] ), .IN4(n6145), 
        .Q(n3684) );
  AO22X1 U4715 ( .IN1(n6886), .IN2(n6142), .IN3(\FIFO[27][18] ), .IN4(n6145), 
        .Q(n3685) );
  AO22X1 U4716 ( .IN1(n6875), .IN2(n6141), .IN3(\FIFO[27][19] ), .IN4(n6145), 
        .Q(n3686) );
  AO22X1 U4717 ( .IN1(n6853), .IN2(n6141), .IN3(\FIFO[27][21] ), .IN4(n6145), 
        .Q(n3688) );
  AO22X1 U4718 ( .IN1(n6842), .IN2(n6141), .IN3(\FIFO[27][22] ), .IN4(n6145), 
        .Q(n3689) );
  AO22X1 U4719 ( .IN1(n6831), .IN2(n6141), .IN3(\FIFO[27][23] ), .IN4(n6145), 
        .Q(n3690) );
  AO22X1 U4720 ( .IN1(n7090), .IN2(n6137), .IN3(\FIFO[26][0] ), .IN4(n6138), 
        .Q(n3699) );
  AO22X1 U4721 ( .IN1(n7073), .IN2(n6136), .IN3(\FIFO[26][1] ), .IN4(n6138), 
        .Q(n3700) );
  AO22X1 U4722 ( .IN1(n7062), .IN2(n6135), .IN3(\FIFO[26][2] ), .IN4(n6138), 
        .Q(n3701) );
  AO22X1 U4723 ( .IN1(n7051), .IN2(n6137), .IN3(\FIFO[26][3] ), .IN4(n6138), 
        .Q(n3702) );
  AO22X1 U4724 ( .IN1(n7040), .IN2(n6136), .IN3(\FIFO[26][4] ), .IN4(n6138), 
        .Q(n3703) );
  AO22X1 U4725 ( .IN1(n7018), .IN2(n6137), .IN3(\FIFO[26][6] ), .IN4(n6138), 
        .Q(n3705) );
  AO22X1 U4726 ( .IN1(n7007), .IN2(n6137), .IN3(\FIFO[26][7] ), .IN4(n6138), 
        .Q(n3706) );
  AO22X1 U4727 ( .IN1(n6996), .IN2(n6137), .IN3(\FIFO[26][8] ), .IN4(n6138), 
        .Q(n3707) );
  AO22X1 U4728 ( .IN1(n6985), .IN2(n6137), .IN3(\FIFO[26][9] ), .IN4(n6138), 
        .Q(n3708) );
  AO22X1 U4729 ( .IN1(n6974), .IN2(n6137), .IN3(\FIFO[26][10] ), .IN4(n6138), 
        .Q(n3709) );
  AO22X1 U4730 ( .IN1(n6963), .IN2(n6137), .IN3(\FIFO[26][11] ), .IN4(n6138), 
        .Q(n3710) );
  AO22X1 U4731 ( .IN1(n6952), .IN2(n6137), .IN3(\FIFO[26][12] ), .IN4(n6139), 
        .Q(n3711) );
  AO22X1 U4732 ( .IN1(n6941), .IN2(n6137), .IN3(\FIFO[26][13] ), .IN4(n6139), 
        .Q(n3712) );
  AO22X1 U4733 ( .IN1(n6930), .IN2(n6136), .IN3(\FIFO[26][14] ), .IN4(n6139), 
        .Q(n3713) );
  AO22X1 U4734 ( .IN1(n6919), .IN2(n6136), .IN3(\FIFO[26][15] ), .IN4(n6139), 
        .Q(n3714) );
  AO22X1 U4735 ( .IN1(n6908), .IN2(n6136), .IN3(\FIFO[26][16] ), .IN4(n6139), 
        .Q(n3715) );
  AO22X1 U4736 ( .IN1(n6897), .IN2(n6136), .IN3(\FIFO[26][17] ), .IN4(n6139), 
        .Q(n3716) );
  AO22X1 U4737 ( .IN1(n6886), .IN2(n6136), .IN3(\FIFO[26][18] ), .IN4(n6139), 
        .Q(n3717) );
  AO22X1 U4738 ( .IN1(n6875), .IN2(n6136), .IN3(\FIFO[26][19] ), .IN4(n6139), 
        .Q(n3718) );
  AO22X1 U4739 ( .IN1(n6864), .IN2(n6136), .IN3(\FIFO[26][20] ), .IN4(n6139), 
        .Q(n3719) );
  AO22X1 U4740 ( .IN1(n6842), .IN2(n6135), .IN3(\FIFO[26][22] ), .IN4(n6139), 
        .Q(n3721) );
  AO22X1 U4741 ( .IN1(n6831), .IN2(n6135), .IN3(\FIFO[26][23] ), .IN4(n6139), 
        .Q(n3722) );
  AO22X1 U4742 ( .IN1(n7089), .IN2(n6119), .IN3(\FIFO[23][0] ), .IN4(n6120), 
        .Q(n3795) );
  AO22X1 U4743 ( .IN1(n7072), .IN2(n6119), .IN3(\FIFO[23][1] ), .IN4(n6120), 
        .Q(n3796) );
  AO22X1 U4744 ( .IN1(n7061), .IN2(n6119), .IN3(\FIFO[23][2] ), .IN4(n6120), 
        .Q(n3797) );
  AO22X1 U4745 ( .IN1(n7050), .IN2(n6119), .IN3(\FIFO[23][3] ), .IN4(n6120), 
        .Q(n3798) );
  AO22X1 U4746 ( .IN1(n7039), .IN2(n6119), .IN3(\FIFO[23][4] ), .IN4(n6120), 
        .Q(n3799) );
  AO22X1 U4747 ( .IN1(n7028), .IN2(n6119), .IN3(\FIFO[23][5] ), .IN4(n6120), 
        .Q(n3800) );
  AO22X1 U4748 ( .IN1(n7017), .IN2(n6119), .IN3(\FIFO[23][6] ), .IN4(n6120), 
        .Q(n3801) );
  AO22X1 U4749 ( .IN1(n7006), .IN2(n6118), .IN3(\FIFO[23][7] ), .IN4(n6120), 
        .Q(n3802) );
  AO22X1 U4750 ( .IN1(n6984), .IN2(n6118), .IN3(\FIFO[23][9] ), .IN4(n6120), 
        .Q(n3804) );
  AO22X1 U4751 ( .IN1(n6973), .IN2(n6118), .IN3(\FIFO[23][10] ), .IN4(n6120), 
        .Q(n3805) );
  AO22X1 U4752 ( .IN1(n6962), .IN2(n6118), .IN3(\FIFO[23][11] ), .IN4(n6120), 
        .Q(n3806) );
  AO22X1 U4753 ( .IN1(n6951), .IN2(n6118), .IN3(\FIFO[23][12] ), .IN4(n6121), 
        .Q(n3807) );
  AO22X1 U4754 ( .IN1(n6940), .IN2(n6118), .IN3(\FIFO[23][13] ), .IN4(n6121), 
        .Q(n3808) );
  AO22X1 U4755 ( .IN1(n6929), .IN2(n6117), .IN3(\FIFO[23][14] ), .IN4(n6121), 
        .Q(n3809) );
  AO22X1 U4756 ( .IN1(n6918), .IN2(n6117), .IN3(\FIFO[23][15] ), .IN4(n6121), 
        .Q(n3810) );
  AO22X1 U4757 ( .IN1(n6907), .IN2(n6117), .IN3(\FIFO[23][16] ), .IN4(n6121), 
        .Q(n3811) );
  AO22X1 U4758 ( .IN1(n6896), .IN2(n6117), .IN3(\FIFO[23][17] ), .IN4(n6121), 
        .Q(n3812) );
  AO22X1 U4759 ( .IN1(n6885), .IN2(n6117), .IN3(\FIFO[23][18] ), .IN4(n6121), 
        .Q(n3813) );
  AO22X1 U4760 ( .IN1(n6874), .IN2(n6117), .IN3(\FIFO[23][19] ), .IN4(n6121), 
        .Q(n3814) );
  AO22X1 U4761 ( .IN1(n6863), .IN2(n6117), .IN3(\FIFO[23][20] ), .IN4(n6121), 
        .Q(n3815) );
  AO22X1 U4762 ( .IN1(n6852), .IN2(n6119), .IN3(\FIFO[23][21] ), .IN4(n6121), 
        .Q(n3816) );
  AO22X1 U4763 ( .IN1(n6841), .IN2(n6118), .IN3(\FIFO[23][22] ), .IN4(n6121), 
        .Q(n3817) );
  AO22X1 U4764 ( .IN1(n6830), .IN2(n6117), .IN3(\FIFO[23][23] ), .IN4(n6121), 
        .Q(n3818) );
  AO22X1 U4765 ( .IN1(n7089), .IN2(n6113), .IN3(\FIFO[22][0] ), .IN4(n6114), 
        .Q(n3827) );
  AO22X1 U4766 ( .IN1(n7072), .IN2(n6113), .IN3(\FIFO[22][1] ), .IN4(n6114), 
        .Q(n3828) );
  AO22X1 U4767 ( .IN1(n7061), .IN2(n6113), .IN3(\FIFO[22][2] ), .IN4(n6114), 
        .Q(n3829) );
  AO22X1 U4768 ( .IN1(n7050), .IN2(n6113), .IN3(\FIFO[22][3] ), .IN4(n6114), 
        .Q(n3830) );
  AO22X1 U4769 ( .IN1(n7039), .IN2(n6113), .IN3(\FIFO[22][4] ), .IN4(n6114), 
        .Q(n3831) );
  AO22X1 U4770 ( .IN1(n7028), .IN2(n6113), .IN3(\FIFO[22][5] ), .IN4(n6114), 
        .Q(n3832) );
  AO22X1 U4771 ( .IN1(n7017), .IN2(n6113), .IN3(\FIFO[22][6] ), .IN4(n6114), 
        .Q(n3833) );
  AO22X1 U4772 ( .IN1(n7006), .IN2(n6112), .IN3(\FIFO[22][7] ), .IN4(n6114), 
        .Q(n3834) );
  AO22X1 U4773 ( .IN1(n6995), .IN2(n6112), .IN3(\FIFO[22][8] ), .IN4(n6114), 
        .Q(n3835) );
  AO22X1 U4774 ( .IN1(n6973), .IN2(n6112), .IN3(\FIFO[22][10] ), .IN4(n6114), 
        .Q(n3837) );
  AO22X1 U4775 ( .IN1(n6962), .IN2(n6112), .IN3(\FIFO[22][11] ), .IN4(n6114), 
        .Q(n3838) );
  AO22X1 U4776 ( .IN1(n6951), .IN2(n6112), .IN3(\FIFO[22][12] ), .IN4(n6115), 
        .Q(n3839) );
  AO22X1 U4777 ( .IN1(n6940), .IN2(n6112), .IN3(\FIFO[22][13] ), .IN4(n6115), 
        .Q(n3840) );
  AO22X1 U4778 ( .IN1(n6929), .IN2(n6113), .IN3(\FIFO[22][14] ), .IN4(n6115), 
        .Q(n3841) );
  AO22X1 U4779 ( .IN1(n6918), .IN2(n6112), .IN3(\FIFO[22][15] ), .IN4(n6115), 
        .Q(n3842) );
  AO22X1 U4780 ( .IN1(n6907), .IN2(n6111), .IN3(\FIFO[22][16] ), .IN4(n6115), 
        .Q(n3843) );
  AO22X1 U4781 ( .IN1(n6896), .IN2(n6113), .IN3(\FIFO[22][17] ), .IN4(n6115), 
        .Q(n3844) );
  AO22X1 U4782 ( .IN1(n6885), .IN2(n6112), .IN3(\FIFO[22][18] ), .IN4(n6115), 
        .Q(n3845) );
  AO22X1 U4783 ( .IN1(n6874), .IN2(n6111), .IN3(\FIFO[22][19] ), .IN4(n6115), 
        .Q(n3846) );
  AO22X1 U4784 ( .IN1(n6863), .IN2(n6113), .IN3(\FIFO[22][20] ), .IN4(n6115), 
        .Q(n3847) );
  AO22X1 U4785 ( .IN1(n6852), .IN2(n6111), .IN3(\FIFO[22][21] ), .IN4(n6115), 
        .Q(n3848) );
  AO22X1 U4786 ( .IN1(n6830), .IN2(n6111), .IN3(\FIFO[22][23] ), .IN4(n6115), 
        .Q(n3850) );
  AO22X1 U4787 ( .IN1(n7072), .IN2(n6095), .IN3(\FIFO[19][1] ), .IN4(n6096), 
        .Q(n3924) );
  AO22X1 U4788 ( .IN1(n7061), .IN2(n6095), .IN3(\FIFO[19][2] ), .IN4(n6096), 
        .Q(n3925) );
  AO22X1 U4789 ( .IN1(n7050), .IN2(n6095), .IN3(\FIFO[19][3] ), .IN4(n6096), 
        .Q(n3926) );
  AO22X1 U4790 ( .IN1(n7039), .IN2(n6095), .IN3(\FIFO[19][4] ), .IN4(n6096), 
        .Q(n3927) );
  AO22X1 U4791 ( .IN1(n7028), .IN2(n6095), .IN3(\FIFO[19][5] ), .IN4(n6096), 
        .Q(n3928) );
  AO22X1 U4792 ( .IN1(n7017), .IN2(n6095), .IN3(\FIFO[19][6] ), .IN4(n6096), 
        .Q(n3929) );
  AO22X1 U4793 ( .IN1(n7006), .IN2(n6094), .IN3(\FIFO[19][7] ), .IN4(n6096), 
        .Q(n3930) );
  AO22X1 U4794 ( .IN1(n6995), .IN2(n6094), .IN3(\FIFO[19][8] ), .IN4(n6096), 
        .Q(n3931) );
  AO22X1 U4795 ( .IN1(n6984), .IN2(n6094), .IN3(\FIFO[19][9] ), .IN4(n6096), 
        .Q(n3932) );
  AO22X1 U4796 ( .IN1(n6973), .IN2(n6094), .IN3(\FIFO[19][10] ), .IN4(n6096), 
        .Q(n3933) );
  AO22X1 U4797 ( .IN1(n6962), .IN2(n6094), .IN3(\FIFO[19][11] ), .IN4(n6096), 
        .Q(n3934) );
  AO22X1 U4798 ( .IN1(n6940), .IN2(n6094), .IN3(\FIFO[19][13] ), .IN4(n6097), 
        .Q(n3936) );
  AO22X1 U4799 ( .IN1(n6929), .IN2(n6093), .IN3(\FIFO[19][14] ), .IN4(n6097), 
        .Q(n3937) );
  AO22X1 U4800 ( .IN1(n6918), .IN2(n6093), .IN3(\FIFO[19][15] ), .IN4(n6097), 
        .Q(n3938) );
  AO22X1 U4801 ( .IN1(n6907), .IN2(n6093), .IN3(\FIFO[19][16] ), .IN4(n6097), 
        .Q(n3939) );
  AO22X1 U4802 ( .IN1(n6896), .IN2(n6093), .IN3(\FIFO[19][17] ), .IN4(n6097), 
        .Q(n3940) );
  AO22X1 U4803 ( .IN1(n6885), .IN2(n6093), .IN3(\FIFO[19][18] ), .IN4(n6097), 
        .Q(n3941) );
  AO22X1 U4804 ( .IN1(n6874), .IN2(n6093), .IN3(\FIFO[19][19] ), .IN4(n6097), 
        .Q(n3942) );
  AO22X1 U4805 ( .IN1(n6863), .IN2(n6093), .IN3(\FIFO[19][20] ), .IN4(n6097), 
        .Q(n3943) );
  AO22X1 U4806 ( .IN1(n6852), .IN2(n6095), .IN3(\FIFO[19][21] ), .IN4(n6097), 
        .Q(n3944) );
  AO22X1 U4807 ( .IN1(n6841), .IN2(n6094), .IN3(\FIFO[19][22] ), .IN4(n6097), 
        .Q(n3945) );
  AO22X1 U4808 ( .IN1(n6830), .IN2(n6093), .IN3(\FIFO[19][23] ), .IN4(n6097), 
        .Q(n3946) );
  AO22X1 U4809 ( .IN1(n7089), .IN2(n6089), .IN3(\FIFO[18][0] ), .IN4(n6090), 
        .Q(n3955) );
  AO22X1 U4810 ( .IN1(n7061), .IN2(n6089), .IN3(\FIFO[18][2] ), .IN4(n6090), 
        .Q(n3957) );
  AO22X1 U4811 ( .IN1(n7050), .IN2(n6089), .IN3(\FIFO[18][3] ), .IN4(n6090), 
        .Q(n3958) );
  AO22X1 U4812 ( .IN1(n7039), .IN2(n6089), .IN3(\FIFO[18][4] ), .IN4(n6090), 
        .Q(n3959) );
  AO22X1 U4813 ( .IN1(n7028), .IN2(n6089), .IN3(\FIFO[18][5] ), .IN4(n6090), 
        .Q(n3960) );
  AO22X1 U4814 ( .IN1(n7017), .IN2(n6089), .IN3(\FIFO[18][6] ), .IN4(n6090), 
        .Q(n3961) );
  AO22X1 U4815 ( .IN1(n7006), .IN2(n6088), .IN3(\FIFO[18][7] ), .IN4(n6090), 
        .Q(n3962) );
  AO22X1 U4816 ( .IN1(n6995), .IN2(n6088), .IN3(\FIFO[18][8] ), .IN4(n6090), 
        .Q(n3963) );
  AO22X1 U4817 ( .IN1(n6984), .IN2(n6088), .IN3(\FIFO[18][9] ), .IN4(n6090), 
        .Q(n3964) );
  AO22X1 U4818 ( .IN1(n6973), .IN2(n6088), .IN3(\FIFO[18][10] ), .IN4(n6090), 
        .Q(n3965) );
  AO22X1 U4819 ( .IN1(n6962), .IN2(n6088), .IN3(\FIFO[18][11] ), .IN4(n6090), 
        .Q(n3966) );
  AO22X1 U4820 ( .IN1(n6951), .IN2(n6088), .IN3(\FIFO[18][12] ), .IN4(n6091), 
        .Q(n3967) );
  AO22X1 U4821 ( .IN1(n6929), .IN2(n6087), .IN3(\FIFO[18][14] ), .IN4(n6091), 
        .Q(n3969) );
  AO22X1 U4822 ( .IN1(n6918), .IN2(n6087), .IN3(\FIFO[18][15] ), .IN4(n6091), 
        .Q(n3970) );
  AO22X1 U4823 ( .IN1(n6907), .IN2(n6087), .IN3(\FIFO[18][16] ), .IN4(n6091), 
        .Q(n3971) );
  AO22X1 U4824 ( .IN1(n6896), .IN2(n6087), .IN3(\FIFO[18][17] ), .IN4(n6091), 
        .Q(n3972) );
  AO22X1 U4825 ( .IN1(n6885), .IN2(n6087), .IN3(\FIFO[18][18] ), .IN4(n6091), 
        .Q(n3973) );
  AO22X1 U4826 ( .IN1(n6874), .IN2(n6087), .IN3(\FIFO[18][19] ), .IN4(n6091), 
        .Q(n3974) );
  AO22X1 U4827 ( .IN1(n6863), .IN2(n6087), .IN3(\FIFO[18][20] ), .IN4(n6091), 
        .Q(n3975) );
  AO22X1 U4828 ( .IN1(n6852), .IN2(n6089), .IN3(\FIFO[18][21] ), .IN4(n6091), 
        .Q(n3976) );
  AO22X1 U4829 ( .IN1(n6841), .IN2(n6088), .IN3(\FIFO[18][22] ), .IN4(n6091), 
        .Q(n3977) );
  AO22X1 U4830 ( .IN1(n6830), .IN2(n6087), .IN3(\FIFO[18][23] ), .IN4(n6091), 
        .Q(n3978) );
  AO22X1 U4831 ( .IN1(n7089), .IN2(n6071), .IN3(\FIFO[15][0] ), .IN4(n6072), 
        .Q(n4051) );
  AO22X1 U4832 ( .IN1(n7072), .IN2(n6071), .IN3(\FIFO[15][1] ), .IN4(n6072), 
        .Q(n4052) );
  AO22X1 U4833 ( .IN1(n7050), .IN2(n6071), .IN3(\FIFO[15][3] ), .IN4(n6072), 
        .Q(n4054) );
  AO22X1 U4834 ( .IN1(n7039), .IN2(n6071), .IN3(\FIFO[15][4] ), .IN4(n6072), 
        .Q(n4055) );
  AO22X1 U4835 ( .IN1(n7028), .IN2(n6071), .IN3(\FIFO[15][5] ), .IN4(n6072), 
        .Q(n4056) );
  AO22X1 U4836 ( .IN1(n7017), .IN2(n6071), .IN3(\FIFO[15][6] ), .IN4(n6072), 
        .Q(n4057) );
  AO22X1 U4837 ( .IN1(n7006), .IN2(n6070), .IN3(\FIFO[15][7] ), .IN4(n6072), 
        .Q(n4058) );
  AO22X1 U4838 ( .IN1(n6995), .IN2(n6070), .IN3(\FIFO[15][8] ), .IN4(n6072), 
        .Q(n4059) );
  AO22X1 U4839 ( .IN1(n6984), .IN2(n6070), .IN3(\FIFO[15][9] ), .IN4(n6072), 
        .Q(n4060) );
  AO22X1 U4840 ( .IN1(n6973), .IN2(n6070), .IN3(\FIFO[15][10] ), .IN4(n6072), 
        .Q(n4061) );
  AO22X1 U4841 ( .IN1(n6962), .IN2(n6070), .IN3(\FIFO[15][11] ), .IN4(n6072), 
        .Q(n4062) );
  AO22X1 U4842 ( .IN1(n6951), .IN2(n6070), .IN3(\FIFO[15][12] ), .IN4(n6073), 
        .Q(n4063) );
  AO22X1 U4843 ( .IN1(n6940), .IN2(n6070), .IN3(\FIFO[15][13] ), .IN4(n6073), 
        .Q(n4064) );
  AO22X1 U4844 ( .IN1(n6918), .IN2(n6069), .IN3(\FIFO[15][15] ), .IN4(n6073), 
        .Q(n4066) );
  AO22X1 U4845 ( .IN1(n6907), .IN2(n6069), .IN3(\FIFO[15][16] ), .IN4(n6073), 
        .Q(n4067) );
  AO22X1 U4846 ( .IN1(n6896), .IN2(n6069), .IN3(\FIFO[15][17] ), .IN4(n6073), 
        .Q(n4068) );
  AO22X1 U4847 ( .IN1(n6885), .IN2(n6069), .IN3(\FIFO[15][18] ), .IN4(n6073), 
        .Q(n4069) );
  AO22X1 U4848 ( .IN1(n6874), .IN2(n6069), .IN3(\FIFO[15][19] ), .IN4(n6073), 
        .Q(n4070) );
  AO22X1 U4849 ( .IN1(n6863), .IN2(n6069), .IN3(\FIFO[15][20] ), .IN4(n6073), 
        .Q(n4071) );
  AO22X1 U4850 ( .IN1(n6852), .IN2(n6071), .IN3(\FIFO[15][21] ), .IN4(n6073), 
        .Q(n4072) );
  AO22X1 U4851 ( .IN1(n6841), .IN2(n6070), .IN3(\FIFO[15][22] ), .IN4(n6073), 
        .Q(n4073) );
  AO22X1 U4852 ( .IN1(n6830), .IN2(n6069), .IN3(\FIFO[15][23] ), .IN4(n6073), 
        .Q(n4074) );
  AO22X1 U4853 ( .IN1(n7089), .IN2(n6065), .IN3(\FIFO[14][0] ), .IN4(n6066), 
        .Q(n4083) );
  AO22X1 U4854 ( .IN1(n7072), .IN2(n6065), .IN3(\FIFO[14][1] ), .IN4(n6066), 
        .Q(n4084) );
  AO22X1 U4855 ( .IN1(n7061), .IN2(n6065), .IN3(\FIFO[14][2] ), .IN4(n6066), 
        .Q(n4085) );
  AO22X1 U4856 ( .IN1(n7039), .IN2(n6065), .IN3(\FIFO[14][4] ), .IN4(n6066), 
        .Q(n4087) );
  AO22X1 U4857 ( .IN1(n7028), .IN2(n6065), .IN3(\FIFO[14][5] ), .IN4(n6066), 
        .Q(n4088) );
  AO22X1 U4858 ( .IN1(n7017), .IN2(n6065), .IN3(\FIFO[14][6] ), .IN4(n6066), 
        .Q(n4089) );
  AO22X1 U4859 ( .IN1(n7006), .IN2(n6064), .IN3(\FIFO[14][7] ), .IN4(n6066), 
        .Q(n4090) );
  AO22X1 U4860 ( .IN1(n6995), .IN2(n6064), .IN3(\FIFO[14][8] ), .IN4(n6066), 
        .Q(n4091) );
  AO22X1 U4861 ( .IN1(n6984), .IN2(n6064), .IN3(\FIFO[14][9] ), .IN4(n6066), 
        .Q(n4092) );
  AO22X1 U4862 ( .IN1(n6973), .IN2(n6064), .IN3(\FIFO[14][10] ), .IN4(n6066), 
        .Q(n4093) );
  AO22X1 U4863 ( .IN1(n6962), .IN2(n6064), .IN3(\FIFO[14][11] ), .IN4(n6066), 
        .Q(n4094) );
  AO22X1 U4864 ( .IN1(n6951), .IN2(n6064), .IN3(\FIFO[14][12] ), .IN4(n6067), 
        .Q(n4095) );
  AO22X1 U4865 ( .IN1(n6940), .IN2(n6064), .IN3(\FIFO[14][13] ), .IN4(n6067), 
        .Q(n4096) );
  AO22X1 U4866 ( .IN1(n6929), .IN2(n6063), .IN3(\FIFO[14][14] ), .IN4(n6067), 
        .Q(n4097) );
  AO22X1 U4867 ( .IN1(n6907), .IN2(n6063), .IN3(\FIFO[14][16] ), .IN4(n6067), 
        .Q(n4099) );
  AO22X1 U4868 ( .IN1(n6896), .IN2(n6063), .IN3(\FIFO[14][17] ), .IN4(n6067), 
        .Q(n4100) );
  AO22X1 U4869 ( .IN1(n6885), .IN2(n6063), .IN3(\FIFO[14][18] ), .IN4(n6067), 
        .Q(n4101) );
  AO22X1 U4870 ( .IN1(n6874), .IN2(n6063), .IN3(\FIFO[14][19] ), .IN4(n6067), 
        .Q(n4102) );
  AO22X1 U4871 ( .IN1(n6863), .IN2(n6063), .IN3(\FIFO[14][20] ), .IN4(n6067), 
        .Q(n4103) );
  AO22X1 U4872 ( .IN1(n6852), .IN2(n6065), .IN3(\FIFO[14][21] ), .IN4(n6067), 
        .Q(n4104) );
  AO22X1 U4873 ( .IN1(n6841), .IN2(n6064), .IN3(\FIFO[14][22] ), .IN4(n6067), 
        .Q(n4105) );
  AO22X1 U4874 ( .IN1(n6830), .IN2(n6063), .IN3(\FIFO[14][23] ), .IN4(n6067), 
        .Q(n4106) );
  AO22X1 U4875 ( .IN1(n7088), .IN2(n6047), .IN3(\FIFO[11][0] ), .IN4(n6048), 
        .Q(n4179) );
  AO22X1 U4876 ( .IN1(n7071), .IN2(n6047), .IN3(\FIFO[11][1] ), .IN4(n6048), 
        .Q(n4180) );
  AO22X1 U4877 ( .IN1(n7060), .IN2(n6047), .IN3(\FIFO[11][2] ), .IN4(n6048), 
        .Q(n4181) );
  AO22X1 U4878 ( .IN1(n7049), .IN2(n6047), .IN3(\FIFO[11][3] ), .IN4(n6048), 
        .Q(n4182) );
  AO22X1 U4879 ( .IN1(n7027), .IN2(n6047), .IN3(\FIFO[11][5] ), .IN4(n6048), 
        .Q(n4184) );
  AO22X1 U4880 ( .IN1(n7016), .IN2(n6047), .IN3(\FIFO[11][6] ), .IN4(n6048), 
        .Q(n4185) );
  AO22X1 U4881 ( .IN1(n7005), .IN2(n6046), .IN3(\FIFO[11][7] ), .IN4(n6048), 
        .Q(n4186) );
  AO22X1 U4882 ( .IN1(n6994), .IN2(n6046), .IN3(\FIFO[11][8] ), .IN4(n6048), 
        .Q(n4187) );
  AO22X1 U4883 ( .IN1(n6983), .IN2(n6046), .IN3(\FIFO[11][9] ), .IN4(n6048), 
        .Q(n4188) );
  AO22X1 U4884 ( .IN1(n6972), .IN2(n6046), .IN3(\FIFO[11][10] ), .IN4(n6048), 
        .Q(n4189) );
  AO22X1 U4885 ( .IN1(n6961), .IN2(n6046), .IN3(\FIFO[11][11] ), .IN4(n6048), 
        .Q(n4190) );
  AO22X1 U4886 ( .IN1(n6950), .IN2(n6046), .IN3(\FIFO[11][12] ), .IN4(n6049), 
        .Q(n4191) );
  AO22X1 U4887 ( .IN1(n6939), .IN2(n6046), .IN3(\FIFO[11][13] ), .IN4(n6049), 
        .Q(n4192) );
  AO22X1 U4888 ( .IN1(n6928), .IN2(n6045), .IN3(\FIFO[11][14] ), .IN4(n6049), 
        .Q(n4193) );
  AO22X1 U4889 ( .IN1(n6917), .IN2(n6045), .IN3(\FIFO[11][15] ), .IN4(n6049), 
        .Q(n4194) );
  AO22X1 U4890 ( .IN1(n6895), .IN2(n6045), .IN3(\FIFO[11][17] ), .IN4(n6049), 
        .Q(n4196) );
  AO22X1 U4891 ( .IN1(n6884), .IN2(n6045), .IN3(\FIFO[11][18] ), .IN4(n6049), 
        .Q(n4197) );
  AO22X1 U4892 ( .IN1(n6873), .IN2(n6045), .IN3(\FIFO[11][19] ), .IN4(n6049), 
        .Q(n4198) );
  AO22X1 U4893 ( .IN1(n6862), .IN2(n6045), .IN3(\FIFO[11][20] ), .IN4(n6049), 
        .Q(n4199) );
  AO22X1 U4894 ( .IN1(n6851), .IN2(n6047), .IN3(\FIFO[11][21] ), .IN4(n6049), 
        .Q(n4200) );
  AO22X1 U4895 ( .IN1(n6840), .IN2(n6046), .IN3(\FIFO[11][22] ), .IN4(n6049), 
        .Q(n4201) );
  AO22X1 U4896 ( .IN1(n6829), .IN2(n6045), .IN3(\FIFO[11][23] ), .IN4(n6049), 
        .Q(n4202) );
  AO22X1 U4897 ( .IN1(n7088), .IN2(n6041), .IN3(\FIFO[10][0] ), .IN4(n6042), 
        .Q(n4211) );
  AO22X1 U4898 ( .IN1(n7071), .IN2(n6041), .IN3(\FIFO[10][1] ), .IN4(n6042), 
        .Q(n4212) );
  AO22X1 U4899 ( .IN1(n7060), .IN2(n6041), .IN3(\FIFO[10][2] ), .IN4(n6042), 
        .Q(n4213) );
  AO22X1 U4900 ( .IN1(n7049), .IN2(n6041), .IN3(\FIFO[10][3] ), .IN4(n6042), 
        .Q(n4214) );
  AO22X1 U4901 ( .IN1(n7038), .IN2(n6041), .IN3(\FIFO[10][4] ), .IN4(n6042), 
        .Q(n4215) );
  AO22X1 U4902 ( .IN1(n7016), .IN2(n6041), .IN3(\FIFO[10][6] ), .IN4(n6042), 
        .Q(n4217) );
  AO22X1 U4903 ( .IN1(n7005), .IN2(n6040), .IN3(\FIFO[10][7] ), .IN4(n6042), 
        .Q(n4218) );
  AO22X1 U4904 ( .IN1(n6994), .IN2(n6040), .IN3(\FIFO[10][8] ), .IN4(n6042), 
        .Q(n4219) );
  AO22X1 U4905 ( .IN1(n6983), .IN2(n6040), .IN3(\FIFO[10][9] ), .IN4(n6042), 
        .Q(n4220) );
  AO22X1 U4906 ( .IN1(n6972), .IN2(n6040), .IN3(\FIFO[10][10] ), .IN4(n6042), 
        .Q(n4221) );
  AO22X1 U4907 ( .IN1(n6961), .IN2(n6040), .IN3(\FIFO[10][11] ), .IN4(n6042), 
        .Q(n4222) );
  AO22X1 U4908 ( .IN1(n6950), .IN2(n6040), .IN3(\FIFO[10][12] ), .IN4(n6043), 
        .Q(n4223) );
  AO22X1 U4909 ( .IN1(n6939), .IN2(n6040), .IN3(\FIFO[10][13] ), .IN4(n6043), 
        .Q(n4224) );
  AO22X1 U4910 ( .IN1(n6928), .IN2(n6039), .IN3(\FIFO[10][14] ), .IN4(n6043), 
        .Q(n4225) );
  AO22X1 U4911 ( .IN1(n6917), .IN2(n6039), .IN3(\FIFO[10][15] ), .IN4(n6043), 
        .Q(n4226) );
  AO22X1 U4912 ( .IN1(n6906), .IN2(n6039), .IN3(\FIFO[10][16] ), .IN4(n6043), 
        .Q(n4227) );
  AO22X1 U4913 ( .IN1(n6884), .IN2(n6039), .IN3(\FIFO[10][18] ), .IN4(n6043), 
        .Q(n4229) );
  AO22X1 U4914 ( .IN1(n6873), .IN2(n6039), .IN3(\FIFO[10][19] ), .IN4(n6043), 
        .Q(n4230) );
  AO22X1 U4915 ( .IN1(n6862), .IN2(n6039), .IN3(\FIFO[10][20] ), .IN4(n6043), 
        .Q(n4231) );
  AO22X1 U4916 ( .IN1(n6851), .IN2(n6041), .IN3(\FIFO[10][21] ), .IN4(n6043), 
        .Q(n4232) );
  AO22X1 U4917 ( .IN1(n6840), .IN2(n6040), .IN3(\FIFO[10][22] ), .IN4(n6043), 
        .Q(n4233) );
  AO22X1 U4918 ( .IN1(n6829), .IN2(n6039), .IN3(\FIFO[10][23] ), .IN4(n6043), 
        .Q(n4234) );
  AO22X1 U4919 ( .IN1(n7088), .IN2(n6023), .IN3(\FIFO[7][0] ), .IN4(n6024), 
        .Q(n4307) );
  AO22X1 U4920 ( .IN1(n7071), .IN2(n6022), .IN3(\FIFO[7][1] ), .IN4(n6024), 
        .Q(n4308) );
  AO22X1 U4921 ( .IN1(n7049), .IN2(n6023), .IN3(\FIFO[7][3] ), .IN4(n6024), 
        .Q(n4310) );
  AO22X1 U4922 ( .IN1(n7038), .IN2(n6022), .IN3(\FIFO[7][4] ), .IN4(n6024), 
        .Q(n4311) );
  AO22X1 U4923 ( .IN1(n7027), .IN2(n6021), .IN3(\FIFO[7][5] ), .IN4(n6024), 
        .Q(n4312) );
  AO22X1 U4924 ( .IN1(n7016), .IN2(n6023), .IN3(\FIFO[7][6] ), .IN4(n6024), 
        .Q(n4313) );
  AO22X1 U4925 ( .IN1(n7005), .IN2(n6023), .IN3(\FIFO[7][7] ), .IN4(n6024), 
        .Q(n4314) );
  AO22X1 U4926 ( .IN1(n6994), .IN2(n6023), .IN3(\FIFO[7][8] ), .IN4(n6024), 
        .Q(n4315) );
  AO22X1 U4927 ( .IN1(n6983), .IN2(n6023), .IN3(\FIFO[7][9] ), .IN4(n6024), 
        .Q(n4316) );
  AO22X1 U4928 ( .IN1(n6972), .IN2(n6023), .IN3(\FIFO[7][10] ), .IN4(n6024), 
        .Q(n4317) );
  AO22X1 U4929 ( .IN1(n6961), .IN2(n6023), .IN3(\FIFO[7][11] ), .IN4(n6024), 
        .Q(n4318) );
  AO22X1 U4930 ( .IN1(n6950), .IN2(n6023), .IN3(\FIFO[7][12] ), .IN4(n6025), 
        .Q(n4319) );
  AO22X1 U4931 ( .IN1(n6939), .IN2(n6023), .IN3(\FIFO[7][13] ), .IN4(n6025), 
        .Q(n4320) );
  AO22X1 U4932 ( .IN1(n6928), .IN2(n6022), .IN3(\FIFO[7][14] ), .IN4(n6025), 
        .Q(n4321) );
  AO22X1 U4933 ( .IN1(n6917), .IN2(n6022), .IN3(\FIFO[7][15] ), .IN4(n6025), 
        .Q(n4322) );
  AO22X1 U4934 ( .IN1(n6906), .IN2(n6022), .IN3(\FIFO[7][16] ), .IN4(n6025), 
        .Q(n4323) );
  AO22X1 U4935 ( .IN1(n6895), .IN2(n6022), .IN3(\FIFO[7][17] ), .IN4(n6025), 
        .Q(n4324) );
  AO22X1 U4936 ( .IN1(n6884), .IN2(n6022), .IN3(\FIFO[7][18] ), .IN4(n6025), 
        .Q(n4325) );
  AO22X1 U4937 ( .IN1(n6873), .IN2(n6022), .IN3(\FIFO[7][19] ), .IN4(n6025), 
        .Q(n4326) );
  AO22X1 U4938 ( .IN1(n6862), .IN2(n6022), .IN3(\FIFO[7][20] ), .IN4(n6025), 
        .Q(n4327) );
  AO22X1 U4939 ( .IN1(n6840), .IN2(n6021), .IN3(\FIFO[7][22] ), .IN4(n6025), 
        .Q(n4329) );
  AO22X1 U4940 ( .IN1(n6829), .IN2(n6021), .IN3(\FIFO[7][23] ), .IN4(n6025), 
        .Q(n4330) );
  AO22X1 U4941 ( .IN1(n7088), .IN2(n6017), .IN3(\FIFO[6][0] ), .IN4(n6018), 
        .Q(n4339) );
  AO22X1 U4942 ( .IN1(n7071), .IN2(n6017), .IN3(\FIFO[6][1] ), .IN4(n6018), 
        .Q(n4340) );
  AO22X1 U4943 ( .IN1(n7060), .IN2(n6017), .IN3(\FIFO[6][2] ), .IN4(n6018), 
        .Q(n4341) );
  AO22X1 U4944 ( .IN1(n7049), .IN2(n6017), .IN3(\FIFO[6][3] ), .IN4(n6018), 
        .Q(n4342) );
  AO22X1 U4945 ( .IN1(n7038), .IN2(n6017), .IN3(\FIFO[6][4] ), .IN4(n6018), 
        .Q(n4343) );
  AO22X1 U4946 ( .IN1(n7027), .IN2(n6017), .IN3(\FIFO[6][5] ), .IN4(n6018), 
        .Q(n4344) );
  AO22X1 U4947 ( .IN1(n7016), .IN2(n6017), .IN3(\FIFO[6][6] ), .IN4(n6018), 
        .Q(n4345) );
  AO22X1 U4948 ( .IN1(n7005), .IN2(n6016), .IN3(\FIFO[6][7] ), .IN4(n6018), 
        .Q(n4346) );
  AO22X1 U4949 ( .IN1(n6983), .IN2(n6016), .IN3(\FIFO[6][9] ), .IN4(n6018), 
        .Q(n4348) );
  AO22X1 U4950 ( .IN1(n6972), .IN2(n6016), .IN3(\FIFO[6][10] ), .IN4(n6018), 
        .Q(n4349) );
  AO22X1 U4951 ( .IN1(n6961), .IN2(n6016), .IN3(\FIFO[6][11] ), .IN4(n6018), 
        .Q(n4350) );
  AO22X1 U4952 ( .IN1(n6950), .IN2(n6016), .IN3(\FIFO[6][12] ), .IN4(n6019), 
        .Q(n4351) );
  AO22X1 U4953 ( .IN1(n6939), .IN2(n6016), .IN3(\FIFO[6][13] ), .IN4(n6019), 
        .Q(n4352) );
  AO22X1 U4954 ( .IN1(n6928), .IN2(n6015), .IN3(\FIFO[6][14] ), .IN4(n6019), 
        .Q(n4353) );
  AO22X1 U4955 ( .IN1(n6917), .IN2(n6015), .IN3(\FIFO[6][15] ), .IN4(n6019), 
        .Q(n4354) );
  AO22X1 U4956 ( .IN1(n6906), .IN2(n6015), .IN3(\FIFO[6][16] ), .IN4(n6019), 
        .Q(n4355) );
  AO22X1 U4957 ( .IN1(n6895), .IN2(n6015), .IN3(\FIFO[6][17] ), .IN4(n6019), 
        .Q(n4356) );
  AO22X1 U4958 ( .IN1(n6884), .IN2(n6015), .IN3(\FIFO[6][18] ), .IN4(n6019), 
        .Q(n4357) );
  AO22X1 U4959 ( .IN1(n6862), .IN2(n6015), .IN3(\FIFO[6][20] ), .IN4(n6019), 
        .Q(n4359) );
  AO22X1 U4960 ( .IN1(n6851), .IN2(n6017), .IN3(\FIFO[6][21] ), .IN4(n6019), 
        .Q(n4360) );
  AO22X1 U4961 ( .IN1(n6840), .IN2(n6016), .IN3(\FIFO[6][22] ), .IN4(n6019), 
        .Q(n4361) );
  AO22X1 U4962 ( .IN1(n6829), .IN2(n6015), .IN3(\FIFO[6][23] ), .IN4(n6019), 
        .Q(n4362) );
  AO22X1 U4963 ( .IN1(n7088), .IN2(n5999), .IN3(\FIFO[3][0] ), .IN4(n6000), 
        .Q(n4435) );
  AO22X1 U4964 ( .IN1(n7071), .IN2(n5999), .IN3(\FIFO[3][1] ), .IN4(n6000), 
        .Q(n4436) );
  AO22X1 U4965 ( .IN1(n7060), .IN2(n5999), .IN3(\FIFO[3][2] ), .IN4(n6000), 
        .Q(n4437) );
  AO22X1 U4966 ( .IN1(n7049), .IN2(n5999), .IN3(\FIFO[3][3] ), .IN4(n6000), 
        .Q(n4438) );
  AO22X1 U4967 ( .IN1(n7038), .IN2(n5999), .IN3(\FIFO[3][4] ), .IN4(n6000), 
        .Q(n4439) );
  AO22X1 U4968 ( .IN1(n7027), .IN2(n5999), .IN3(\FIFO[3][5] ), .IN4(n6000), 
        .Q(n4440) );
  AO22X1 U4969 ( .IN1(n7016), .IN2(n5999), .IN3(\FIFO[3][6] ), .IN4(n6000), 
        .Q(n4441) );
  AO22X1 U4970 ( .IN1(n7005), .IN2(n5998), .IN3(\FIFO[3][7] ), .IN4(n6000), 
        .Q(n4442) );
  AO22X1 U4971 ( .IN1(n6994), .IN2(n5998), .IN3(\FIFO[3][8] ), .IN4(n6000), 
        .Q(n4443) );
  AO22X1 U4972 ( .IN1(n6983), .IN2(n5998), .IN3(\FIFO[3][9] ), .IN4(n6000), 
        .Q(n4444) );
  AO22X1 U4973 ( .IN1(n6972), .IN2(n5998), .IN3(\FIFO[3][10] ), .IN4(n6000), 
        .Q(n4445) );
  AO22X1 U4974 ( .IN1(n6961), .IN2(n5998), .IN3(\FIFO[3][11] ), .IN4(n6000), 
        .Q(n4446) );
  AO22X1 U4975 ( .IN1(n6950), .IN2(n5998), .IN3(\FIFO[3][12] ), .IN4(n6001), 
        .Q(n4447) );
  AO22X1 U4976 ( .IN1(n6939), .IN2(n5998), .IN3(\FIFO[3][13] ), .IN4(n6001), 
        .Q(n4448) );
  AO22X1 U4977 ( .IN1(n6928), .IN2(n5999), .IN3(\FIFO[3][14] ), .IN4(n6001), 
        .Q(n4449) );
  AO22X1 U4978 ( .IN1(n6906), .IN2(n5997), .IN3(\FIFO[3][16] ), .IN4(n6001), 
        .Q(n4451) );
  AO22X1 U4979 ( .IN1(n6895), .IN2(n5999), .IN3(\FIFO[3][17] ), .IN4(n6001), 
        .Q(n4452) );
  AO22X1 U4980 ( .IN1(n6884), .IN2(n5998), .IN3(\FIFO[3][18] ), .IN4(n6001), 
        .Q(n4453) );
  AO22X1 U4981 ( .IN1(n6873), .IN2(n5997), .IN3(\FIFO[3][19] ), .IN4(n6001), 
        .Q(n4454) );
  AO22X1 U4982 ( .IN1(n6862), .IN2(n5999), .IN3(\FIFO[3][20] ), .IN4(n6001), 
        .Q(n4455) );
  AO22X1 U4983 ( .IN1(n6851), .IN2(n5997), .IN3(\FIFO[3][21] ), .IN4(n6001), 
        .Q(n4456) );
  AO22X1 U4984 ( .IN1(n6829), .IN2(n5997), .IN3(\FIFO[3][23] ), .IN4(n6001), 
        .Q(n4458) );
  AO22X1 U4985 ( .IN1(n7088), .IN2(n5993), .IN3(\FIFO[2][0] ), .IN4(n5994), 
        .Q(n4467) );
  AO22X1 U4986 ( .IN1(n7071), .IN2(n5992), .IN3(\FIFO[2][1] ), .IN4(n5994), 
        .Q(n4468) );
  AO22X1 U4987 ( .IN1(n7060), .IN2(n5991), .IN3(\FIFO[2][2] ), .IN4(n5994), 
        .Q(n4469) );
  AO22X1 U4988 ( .IN1(n7038), .IN2(n5992), .IN3(\FIFO[2][4] ), .IN4(n5994), 
        .Q(n4471) );
  AO22X1 U4989 ( .IN1(n7027), .IN2(n5991), .IN3(\FIFO[2][5] ), .IN4(n5994), 
        .Q(n4472) );
  AO22X1 U4990 ( .IN1(n7016), .IN2(n5993), .IN3(\FIFO[2][6] ), .IN4(n5994), 
        .Q(n4473) );
  AO22X1 U4991 ( .IN1(n7005), .IN2(n5993), .IN3(\FIFO[2][7] ), .IN4(n5994), 
        .Q(n4474) );
  AO22X1 U4992 ( .IN1(n6994), .IN2(n5993), .IN3(\FIFO[2][8] ), .IN4(n5994), 
        .Q(n4475) );
  AO22X1 U4993 ( .IN1(n6983), .IN2(n5993), .IN3(\FIFO[2][9] ), .IN4(n5994), 
        .Q(n4476) );
  AO22X1 U4994 ( .IN1(n6972), .IN2(n5993), .IN3(\FIFO[2][10] ), .IN4(n5994), 
        .Q(n4477) );
  AO22X1 U4995 ( .IN1(n6961), .IN2(n5993), .IN3(\FIFO[2][11] ), .IN4(n5994), 
        .Q(n4478) );
  AO22X1 U4996 ( .IN1(n6950), .IN2(n5993), .IN3(\FIFO[2][12] ), .IN4(n5995), 
        .Q(n4479) );
  AO22X1 U4997 ( .IN1(n6939), .IN2(n5993), .IN3(\FIFO[2][13] ), .IN4(n5995), 
        .Q(n4480) );
  AO22X1 U4998 ( .IN1(n6928), .IN2(n5992), .IN3(\FIFO[2][14] ), .IN4(n5995), 
        .Q(n4481) );
  AO22X1 U4999 ( .IN1(n6917), .IN2(n5992), .IN3(\FIFO[2][15] ), .IN4(n5995), 
        .Q(n4482) );
  AO22X1 U5000 ( .IN1(n6906), .IN2(n5992), .IN3(\FIFO[2][16] ), .IN4(n5995), 
        .Q(n4483) );
  AO22X1 U5001 ( .IN1(n6895), .IN2(n5992), .IN3(\FIFO[2][17] ), .IN4(n5995), 
        .Q(n4484) );
  AO22X1 U5002 ( .IN1(n6884), .IN2(n5992), .IN3(\FIFO[2][18] ), .IN4(n5995), 
        .Q(n4485) );
  AO22X1 U5003 ( .IN1(n6873), .IN2(n5992), .IN3(\FIFO[2][19] ), .IN4(n5995), 
        .Q(n4486) );
  AO22X1 U5004 ( .IN1(n6862), .IN2(n5992), .IN3(\FIFO[2][20] ), .IN4(n5995), 
        .Q(n4487) );
  AO22X1 U5005 ( .IN1(n6851), .IN2(n5991), .IN3(\FIFO[2][21] ), .IN4(n5995), 
        .Q(n4488) );
  AO22X1 U5006 ( .IN1(n6840), .IN2(n5991), .IN3(\FIFO[2][22] ), .IN4(n5995), 
        .Q(n4489) );
  AO22X1 U5007 ( .IN1(n7097), .IN2(n6695), .IN3(\FIFO[119][0] ), .IN4(n6696), 
        .Q(n723) );
  AO22X1 U5008 ( .IN1(n7080), .IN2(n6694), .IN3(\FIFO[119][1] ), .IN4(n6696), 
        .Q(n724) );
  AO22X1 U5009 ( .IN1(n7069), .IN2(n6693), .IN3(\FIFO[119][2] ), .IN4(n6696), 
        .Q(n725) );
  AO22X1 U5010 ( .IN1(n7058), .IN2(n6695), .IN3(\FIFO[119][3] ), .IN4(n6696), 
        .Q(n726) );
  AO22X1 U5011 ( .IN1(n7047), .IN2(n6694), .IN3(\FIFO[119][4] ), .IN4(n6696), 
        .Q(n727) );
  AO22X1 U5012 ( .IN1(n7036), .IN2(n6693), .IN3(\FIFO[119][5] ), .IN4(n6696), 
        .Q(n728) );
  AO22X1 U5013 ( .IN1(n7025), .IN2(n6695), .IN3(\FIFO[119][6] ), .IN4(n6696), 
        .Q(n729) );
  AO22X1 U5014 ( .IN1(n7014), .IN2(n6695), .IN3(\FIFO[119][7] ), .IN4(n6696), 
        .Q(n730) );
  AO22X1 U5015 ( .IN1(n7003), .IN2(n6695), .IN3(\FIFO[119][8] ), .IN4(n6696), 
        .Q(n731) );
  AO22X1 U5016 ( .IN1(n6992), .IN2(n6695), .IN3(\FIFO[119][9] ), .IN4(n6696), 
        .Q(n732) );
  AO22X1 U5017 ( .IN1(n6981), .IN2(n6695), .IN3(\FIFO[119][10] ), .IN4(n6696), 
        .Q(n733) );
  AO22X1 U5018 ( .IN1(n6970), .IN2(n6695), .IN3(\FIFO[119][11] ), .IN4(n6696), 
        .Q(n734) );
  AO22X1 U5019 ( .IN1(n6959), .IN2(n6695), .IN3(\FIFO[119][12] ), .IN4(n6697), 
        .Q(n735) );
  AO22X1 U5020 ( .IN1(n6948), .IN2(n6695), .IN3(\FIFO[119][13] ), .IN4(n6697), 
        .Q(n736) );
  AO22X1 U5021 ( .IN1(n6937), .IN2(n6694), .IN3(\FIFO[119][14] ), .IN4(n6697), 
        .Q(n737) );
  AO22X1 U5022 ( .IN1(n6926), .IN2(n6694), .IN3(\FIFO[119][15] ), .IN4(n6697), 
        .Q(n738) );
  AO22X1 U5023 ( .IN1(n6915), .IN2(n6694), .IN3(\FIFO[119][16] ), .IN4(n6697), 
        .Q(n739) );
  AO22X1 U5024 ( .IN1(n6904), .IN2(n6694), .IN3(\FIFO[119][17] ), .IN4(n6697), 
        .Q(n740) );
  AO22X1 U5025 ( .IN1(n6893), .IN2(n6694), .IN3(\FIFO[119][18] ), .IN4(n6697), 
        .Q(n741) );
  AO22X1 U5026 ( .IN1(n6882), .IN2(n6694), .IN3(\FIFO[119][19] ), .IN4(n6697), 
        .Q(n742) );
  AO22X1 U5027 ( .IN1(n6871), .IN2(n6694), .IN3(\FIFO[119][20] ), .IN4(n6697), 
        .Q(n743) );
  AO22X1 U5028 ( .IN1(n6860), .IN2(n6693), .IN3(\FIFO[119][21] ), .IN4(n6697), 
        .Q(n744) );
  AO22X1 U5029 ( .IN1(n6849), .IN2(n6693), .IN3(\FIFO[119][22] ), .IN4(n6697), 
        .Q(n745) );
  AO22X1 U5030 ( .IN1(n6838), .IN2(n6693), .IN3(\FIFO[119][23] ), .IN4(n6697), 
        .Q(n746) );
  AO22X1 U5031 ( .IN1(n7097), .IN2(n6689), .IN3(\FIFO[118][0] ), .IN4(n6690), 
        .Q(n755) );
  AO22X1 U5032 ( .IN1(n7080), .IN2(n6689), .IN3(\FIFO[118][1] ), .IN4(n6690), 
        .Q(n756) );
  AO22X1 U5033 ( .IN1(n7069), .IN2(n6689), .IN3(\FIFO[118][2] ), .IN4(n6690), 
        .Q(n757) );
  AO22X1 U5034 ( .IN1(n7058), .IN2(n6689), .IN3(\FIFO[118][3] ), .IN4(n6690), 
        .Q(n758) );
  AO22X1 U5035 ( .IN1(n7047), .IN2(n6689), .IN3(\FIFO[118][4] ), .IN4(n6690), 
        .Q(n759) );
  AO22X1 U5036 ( .IN1(n7036), .IN2(n6689), .IN3(\FIFO[118][5] ), .IN4(n6690), 
        .Q(n760) );
  AO22X1 U5037 ( .IN1(n7025), .IN2(n6689), .IN3(\FIFO[118][6] ), .IN4(n6690), 
        .Q(n761) );
  AO22X1 U5038 ( .IN1(n7014), .IN2(n6688), .IN3(\FIFO[118][7] ), .IN4(n6690), 
        .Q(n762) );
  AO22X1 U5039 ( .IN1(n7003), .IN2(n6688), .IN3(\FIFO[118][8] ), .IN4(n6690), 
        .Q(n763) );
  AO22X1 U5040 ( .IN1(n6992), .IN2(n6688), .IN3(\FIFO[118][9] ), .IN4(n6690), 
        .Q(n764) );
  AO22X1 U5041 ( .IN1(n6981), .IN2(n6688), .IN3(\FIFO[118][10] ), .IN4(n6690), 
        .Q(n765) );
  AO22X1 U5042 ( .IN1(n6970), .IN2(n6688), .IN3(\FIFO[118][11] ), .IN4(n6690), 
        .Q(n766) );
  AO22X1 U5043 ( .IN1(n6959), .IN2(n6688), .IN3(\FIFO[118][12] ), .IN4(n6691), 
        .Q(n767) );
  AO22X1 U5044 ( .IN1(n6948), .IN2(n6688), .IN3(\FIFO[118][13] ), .IN4(n6691), 
        .Q(n768) );
  AO22X1 U5045 ( .IN1(n6937), .IN2(n6687), .IN3(\FIFO[118][14] ), .IN4(n6691), 
        .Q(n769) );
  AO22X1 U5046 ( .IN1(n6926), .IN2(n6687), .IN3(\FIFO[118][15] ), .IN4(n6691), 
        .Q(n770) );
  AO22X1 U5047 ( .IN1(n6915), .IN2(n6687), .IN3(\FIFO[118][16] ), .IN4(n6691), 
        .Q(n771) );
  AO22X1 U5048 ( .IN1(n6904), .IN2(n6687), .IN3(\FIFO[118][17] ), .IN4(n6691), 
        .Q(n772) );
  AO22X1 U5049 ( .IN1(n6893), .IN2(n6687), .IN3(\FIFO[118][18] ), .IN4(n6691), 
        .Q(n773) );
  AO22X1 U5050 ( .IN1(n6882), .IN2(n6687), .IN3(\FIFO[118][19] ), .IN4(n6691), 
        .Q(n774) );
  AO22X1 U5051 ( .IN1(n6871), .IN2(n6687), .IN3(\FIFO[118][20] ), .IN4(n6691), 
        .Q(n775) );
  AO22X1 U5052 ( .IN1(n6860), .IN2(n256), .IN3(\FIFO[118][21] ), .IN4(n6691), 
        .Q(n776) );
  AO22X1 U5053 ( .IN1(n6849), .IN2(n6689), .IN3(\FIFO[118][22] ), .IN4(n6691), 
        .Q(n777) );
  AO22X1 U5054 ( .IN1(n6838), .IN2(n6688), .IN3(\FIFO[118][23] ), .IN4(n6691), 
        .Q(n778) );
  AO22X1 U5055 ( .IN1(n7097), .IN2(n6671), .IN3(\FIFO[115][0] ), .IN4(n6672), 
        .Q(n851) );
  AO22X1 U5056 ( .IN1(n7080), .IN2(n6671), .IN3(\FIFO[115][1] ), .IN4(n6672), 
        .Q(n852) );
  AO22X1 U5057 ( .IN1(n7069), .IN2(n6671), .IN3(\FIFO[115][2] ), .IN4(n6672), 
        .Q(n853) );
  AO22X1 U5058 ( .IN1(n7058), .IN2(n6671), .IN3(\FIFO[115][3] ), .IN4(n6672), 
        .Q(n854) );
  AO22X1 U5059 ( .IN1(n7047), .IN2(n6671), .IN3(\FIFO[115][4] ), .IN4(n6672), 
        .Q(n855) );
  AO22X1 U5060 ( .IN1(n7036), .IN2(n6671), .IN3(\FIFO[115][5] ), .IN4(n6672), 
        .Q(n856) );
  AO22X1 U5061 ( .IN1(n7014), .IN2(n6670), .IN3(\FIFO[115][7] ), .IN4(n6672), 
        .Q(n858) );
  AO22X1 U5062 ( .IN1(n7003), .IN2(n6670), .IN3(\FIFO[115][8] ), .IN4(n6672), 
        .Q(n859) );
  AO22X1 U5063 ( .IN1(n6992), .IN2(n6670), .IN3(\FIFO[115][9] ), .IN4(n6672), 
        .Q(n860) );
  AO22X1 U5064 ( .IN1(n6981), .IN2(n6670), .IN3(\FIFO[115][10] ), .IN4(n6672), 
        .Q(n861) );
  AO22X1 U5065 ( .IN1(n6970), .IN2(n6670), .IN3(\FIFO[115][11] ), .IN4(n6672), 
        .Q(n862) );
  AO22X1 U5066 ( .IN1(n6959), .IN2(n6670), .IN3(\FIFO[115][12] ), .IN4(n6673), 
        .Q(n863) );
  AO22X1 U5067 ( .IN1(n6948), .IN2(n6670), .IN3(\FIFO[115][13] ), .IN4(n6673), 
        .Q(n864) );
  AO22X1 U5068 ( .IN1(n6937), .IN2(n6671), .IN3(\FIFO[115][14] ), .IN4(n6673), 
        .Q(n865) );
  AO22X1 U5069 ( .IN1(n6926), .IN2(n6670), .IN3(\FIFO[115][15] ), .IN4(n6673), 
        .Q(n866) );
  AO22X1 U5070 ( .IN1(n6915), .IN2(n6669), .IN3(\FIFO[115][16] ), .IN4(n6673), 
        .Q(n867) );
  AO22X1 U5071 ( .IN1(n6904), .IN2(n6671), .IN3(\FIFO[115][17] ), .IN4(n6673), 
        .Q(n868) );
  AO22X1 U5072 ( .IN1(n6893), .IN2(n6670), .IN3(\FIFO[115][18] ), .IN4(n6673), 
        .Q(n869) );
  AO22X1 U5073 ( .IN1(n6882), .IN2(n6669), .IN3(\FIFO[115][19] ), .IN4(n6673), 
        .Q(n870) );
  AO22X1 U5074 ( .IN1(n6871), .IN2(n6671), .IN3(\FIFO[115][20] ), .IN4(n6673), 
        .Q(n871) );
  AO22X1 U5075 ( .IN1(n6860), .IN2(n6669), .IN3(\FIFO[115][21] ), .IN4(n6673), 
        .Q(n872) );
  AO22X1 U5076 ( .IN1(n6849), .IN2(n6669), .IN3(\FIFO[115][22] ), .IN4(n6673), 
        .Q(n873) );
  AO22X1 U5077 ( .IN1(n6838), .IN2(n6669), .IN3(\FIFO[115][23] ), .IN4(n6673), 
        .Q(n874) );
  AO22X1 U5078 ( .IN1(n7097), .IN2(n6665), .IN3(\FIFO[114][0] ), .IN4(n6666), 
        .Q(n883) );
  AO22X1 U5079 ( .IN1(n7080), .IN2(n6664), .IN3(\FIFO[114][1] ), .IN4(n6666), 
        .Q(n884) );
  AO22X1 U5080 ( .IN1(n7069), .IN2(n6663), .IN3(\FIFO[114][2] ), .IN4(n6666), 
        .Q(n885) );
  AO22X1 U5081 ( .IN1(n7058), .IN2(n6665), .IN3(\FIFO[114][3] ), .IN4(n6666), 
        .Q(n886) );
  AO22X1 U5082 ( .IN1(n7047), .IN2(n6664), .IN3(\FIFO[114][4] ), .IN4(n6666), 
        .Q(n887) );
  AO22X1 U5083 ( .IN1(n7036), .IN2(n6663), .IN3(\FIFO[114][5] ), .IN4(n6666), 
        .Q(n888) );
  AO22X1 U5084 ( .IN1(n7025), .IN2(n6665), .IN3(\FIFO[114][6] ), .IN4(n6666), 
        .Q(n889) );
  AO22X1 U5085 ( .IN1(n7014), .IN2(n6665), .IN3(\FIFO[114][7] ), .IN4(n6666), 
        .Q(n890) );
  AO22X1 U5086 ( .IN1(n7003), .IN2(n6665), .IN3(\FIFO[114][8] ), .IN4(n6666), 
        .Q(n891) );
  AO22X1 U5087 ( .IN1(n6992), .IN2(n6665), .IN3(\FIFO[114][9] ), .IN4(n6666), 
        .Q(n892) );
  AO22X1 U5088 ( .IN1(n6981), .IN2(n6665), .IN3(\FIFO[114][10] ), .IN4(n6666), 
        .Q(n893) );
  AO22X1 U5089 ( .IN1(n6970), .IN2(n6665), .IN3(\FIFO[114][11] ), .IN4(n6666), 
        .Q(n894) );
  AO22X1 U5090 ( .IN1(n6959), .IN2(n6665), .IN3(\FIFO[114][12] ), .IN4(n6667), 
        .Q(n895) );
  AO22X1 U5091 ( .IN1(n6948), .IN2(n6665), .IN3(\FIFO[114][13] ), .IN4(n6667), 
        .Q(n896) );
  AO22X1 U5092 ( .IN1(n6937), .IN2(n6664), .IN3(\FIFO[114][14] ), .IN4(n6667), 
        .Q(n897) );
  AO22X1 U5093 ( .IN1(n6926), .IN2(n6664), .IN3(\FIFO[114][15] ), .IN4(n6667), 
        .Q(n898) );
  AO22X1 U5094 ( .IN1(n6915), .IN2(n6664), .IN3(\FIFO[114][16] ), .IN4(n6667), 
        .Q(n899) );
  AO22X1 U5095 ( .IN1(n6904), .IN2(n6664), .IN3(\FIFO[114][17] ), .IN4(n6667), 
        .Q(n900) );
  AO22X1 U5096 ( .IN1(n6893), .IN2(n6664), .IN3(\FIFO[114][18] ), .IN4(n6667), 
        .Q(n901) );
  AO22X1 U5097 ( .IN1(n6882), .IN2(n6664), .IN3(\FIFO[114][19] ), .IN4(n6667), 
        .Q(n902) );
  AO22X1 U5098 ( .IN1(n6871), .IN2(n6664), .IN3(\FIFO[114][20] ), .IN4(n6667), 
        .Q(n903) );
  AO22X1 U5099 ( .IN1(n6860), .IN2(n6663), .IN3(\FIFO[114][21] ), .IN4(n6667), 
        .Q(n904) );
  AO22X1 U5100 ( .IN1(n6849), .IN2(n6663), .IN3(\FIFO[114][22] ), .IN4(n6667), 
        .Q(n905) );
  AO22X1 U5101 ( .IN1(n6838), .IN2(n6663), .IN3(\FIFO[114][23] ), .IN4(n6667), 
        .Q(n906) );
  INVX0 U5102 ( .INP(wraddr[5]), .ZN(n7367) );
  INVX0 U5103 ( .INP(wraddr[6]), .ZN(n7368) );
  AO22X1 U5104 ( .IN1(n7098), .IN2(n7084), .IN3(\FIFO[127][0] ), .IN4(n7085), 
        .Q(n467) );
  AO22X1 U5105 ( .IN1(n7081), .IN2(n7084), .IN3(\FIFO[127][1] ), .IN4(n7085), 
        .Q(n468) );
  AO22X1 U5106 ( .IN1(n7070), .IN2(n7084), .IN3(\FIFO[127][2] ), .IN4(n7085), 
        .Q(n469) );
  AO22X1 U5107 ( .IN1(n7059), .IN2(n7084), .IN3(\FIFO[127][3] ), .IN4(n7085), 
        .Q(n470) );
  AO22X1 U5108 ( .IN1(n7048), .IN2(n7084), .IN3(\FIFO[127][4] ), .IN4(n7085), 
        .Q(n471) );
  AO22X1 U5109 ( .IN1(n7037), .IN2(n7084), .IN3(\FIFO[127][5] ), .IN4(n7085), 
        .Q(n472) );
  AO22X1 U5110 ( .IN1(n7026), .IN2(n7084), .IN3(\FIFO[127][6] ), .IN4(n7085), 
        .Q(n473) );
  AO22X1 U5111 ( .IN1(n7015), .IN2(n7083), .IN3(\FIFO[127][7] ), .IN4(n7085), 
        .Q(n474) );
  AO22X1 U5112 ( .IN1(n7004), .IN2(n7083), .IN3(\FIFO[127][8] ), .IN4(n7085), 
        .Q(n475) );
  AO22X1 U5113 ( .IN1(n6993), .IN2(n7083), .IN3(\FIFO[127][9] ), .IN4(n7085), 
        .Q(n476) );
  AO22X1 U5114 ( .IN1(n6982), .IN2(n7083), .IN3(\FIFO[127][10] ), .IN4(n7085), 
        .Q(n477) );
  AO22X1 U5115 ( .IN1(n6971), .IN2(n7083), .IN3(\FIFO[127][11] ), .IN4(n7085), 
        .Q(n478) );
  AO22X1 U5116 ( .IN1(n6960), .IN2(n7083), .IN3(\FIFO[127][12] ), .IN4(n7086), 
        .Q(n479) );
  AO22X1 U5117 ( .IN1(n6949), .IN2(n7083), .IN3(\FIFO[127][13] ), .IN4(n7086), 
        .Q(n480) );
  AO22X1 U5118 ( .IN1(n6938), .IN2(n7082), .IN3(\FIFO[127][14] ), .IN4(n7086), 
        .Q(n481) );
  AO22X1 U5119 ( .IN1(n6927), .IN2(n7082), .IN3(\FIFO[127][15] ), .IN4(n7086), 
        .Q(n482) );
  AO22X1 U5120 ( .IN1(n6916), .IN2(n7082), .IN3(\FIFO[127][16] ), .IN4(n7086), 
        .Q(n483) );
  AO22X1 U5121 ( .IN1(n6905), .IN2(n7082), .IN3(\FIFO[127][17] ), .IN4(n7086), 
        .Q(n484) );
  AO22X1 U5122 ( .IN1(n6894), .IN2(n7082), .IN3(\FIFO[127][18] ), .IN4(n7086), 
        .Q(n485) );
  AO22X1 U5123 ( .IN1(n6883), .IN2(n7082), .IN3(\FIFO[127][19] ), .IN4(n7086), 
        .Q(n486) );
  AO22X1 U5124 ( .IN1(n6872), .IN2(n7082), .IN3(\FIFO[127][20] ), .IN4(n7086), 
        .Q(n487) );
  AO22X1 U5125 ( .IN1(n6861), .IN2(n7084), .IN3(\FIFO[127][21] ), .IN4(n7086), 
        .Q(n488) );
  AO22X1 U5126 ( .IN1(n6850), .IN2(n7083), .IN3(\FIFO[127][22] ), .IN4(n7086), 
        .Q(n489) );
  AO22X1 U5127 ( .IN1(n6839), .IN2(n7082), .IN3(\FIFO[127][23] ), .IN4(n7086), 
        .Q(n490) );
  AO22X1 U5128 ( .IN1(n7098), .IN2(n6737), .IN3(\FIFO[126][0] ), .IN4(n6738), 
        .Q(n499) );
  AO22X1 U5129 ( .IN1(n7081), .IN2(n6737), .IN3(\FIFO[126][1] ), .IN4(n6738), 
        .Q(n500) );
  AO22X1 U5130 ( .IN1(n7070), .IN2(n6737), .IN3(\FIFO[126][2] ), .IN4(n6738), 
        .Q(n501) );
  AO22X1 U5131 ( .IN1(n7059), .IN2(n6737), .IN3(\FIFO[126][3] ), .IN4(n6738), 
        .Q(n502) );
  AO22X1 U5132 ( .IN1(n7048), .IN2(n6737), .IN3(\FIFO[126][4] ), .IN4(n6738), 
        .Q(n503) );
  AO22X1 U5133 ( .IN1(n7037), .IN2(n6737), .IN3(\FIFO[126][5] ), .IN4(n6738), 
        .Q(n504) );
  AO22X1 U5134 ( .IN1(n7026), .IN2(n6737), .IN3(\FIFO[126][6] ), .IN4(n6738), 
        .Q(n505) );
  AO22X1 U5135 ( .IN1(n7015), .IN2(n6736), .IN3(\FIFO[126][7] ), .IN4(n6738), 
        .Q(n506) );
  AO22X1 U5136 ( .IN1(n7004), .IN2(n6736), .IN3(\FIFO[126][8] ), .IN4(n6738), 
        .Q(n507) );
  AO22X1 U5137 ( .IN1(n6993), .IN2(n6736), .IN3(\FIFO[126][9] ), .IN4(n6738), 
        .Q(n508) );
  AO22X1 U5138 ( .IN1(n6982), .IN2(n6736), .IN3(\FIFO[126][10] ), .IN4(n6738), 
        .Q(n509) );
  AO22X1 U5139 ( .IN1(n6971), .IN2(n6736), .IN3(\FIFO[126][11] ), .IN4(n6738), 
        .Q(n510) );
  AO22X1 U5140 ( .IN1(n6960), .IN2(n6736), .IN3(\FIFO[126][12] ), .IN4(n6739), 
        .Q(n511) );
  AO22X1 U5141 ( .IN1(n6949), .IN2(n6736), .IN3(\FIFO[126][13] ), .IN4(n6739), 
        .Q(n512) );
  AO22X1 U5142 ( .IN1(n6938), .IN2(n6735), .IN3(\FIFO[126][14] ), .IN4(n6739), 
        .Q(n513) );
  AO22X1 U5143 ( .IN1(n6927), .IN2(n6735), .IN3(\FIFO[126][15] ), .IN4(n6739), 
        .Q(n514) );
  AO22X1 U5144 ( .IN1(n6916), .IN2(n6735), .IN3(\FIFO[126][16] ), .IN4(n6739), 
        .Q(n515) );
  AO22X1 U5145 ( .IN1(n6905), .IN2(n6735), .IN3(\FIFO[126][17] ), .IN4(n6739), 
        .Q(n516) );
  AO22X1 U5146 ( .IN1(n6894), .IN2(n6735), .IN3(\FIFO[126][18] ), .IN4(n6739), 
        .Q(n517) );
  AO22X1 U5147 ( .IN1(n6883), .IN2(n6735), .IN3(\FIFO[126][19] ), .IN4(n6739), 
        .Q(n518) );
  AO22X1 U5148 ( .IN1(n6872), .IN2(n6735), .IN3(\FIFO[126][20] ), .IN4(n6739), 
        .Q(n519) );
  AO22X1 U5149 ( .IN1(n6861), .IN2(n6737), .IN3(\FIFO[126][21] ), .IN4(n6739), 
        .Q(n520) );
  AO22X1 U5150 ( .IN1(n6850), .IN2(n6736), .IN3(\FIFO[126][22] ), .IN4(n6739), 
        .Q(n521) );
  AO22X1 U5151 ( .IN1(n6839), .IN2(n6735), .IN3(\FIFO[126][23] ), .IN4(n6739), 
        .Q(n522) );
  AO22X1 U5152 ( .IN1(n7098), .IN2(n6731), .IN3(\FIFO[125][0] ), .IN4(n6732), 
        .Q(n531) );
  AO22X1 U5153 ( .IN1(n7081), .IN2(n6731), .IN3(\FIFO[125][1] ), .IN4(n6732), 
        .Q(n532) );
  AO22X1 U5154 ( .IN1(n7070), .IN2(n6731), .IN3(\FIFO[125][2] ), .IN4(n6732), 
        .Q(n533) );
  AO22X1 U5155 ( .IN1(n7059), .IN2(n6731), .IN3(\FIFO[125][3] ), .IN4(n6732), 
        .Q(n534) );
  AO22X1 U5156 ( .IN1(n7048), .IN2(n6731), .IN3(\FIFO[125][4] ), .IN4(n6732), 
        .Q(n535) );
  AO22X1 U5157 ( .IN1(n7037), .IN2(n6731), .IN3(\FIFO[125][5] ), .IN4(n6732), 
        .Q(n536) );
  AO22X1 U5158 ( .IN1(n7026), .IN2(n6731), .IN3(\FIFO[125][6] ), .IN4(n6732), 
        .Q(n537) );
  AO22X1 U5159 ( .IN1(n7015), .IN2(n6730), .IN3(\FIFO[125][7] ), .IN4(n6732), 
        .Q(n538) );
  AO22X1 U5160 ( .IN1(n7004), .IN2(n6730), .IN3(\FIFO[125][8] ), .IN4(n6732), 
        .Q(n539) );
  AO22X1 U5161 ( .IN1(n6993), .IN2(n6730), .IN3(\FIFO[125][9] ), .IN4(n6732), 
        .Q(n540) );
  AO22X1 U5162 ( .IN1(n6982), .IN2(n6730), .IN3(\FIFO[125][10] ), .IN4(n6732), 
        .Q(n541) );
  AO22X1 U5163 ( .IN1(n6971), .IN2(n6730), .IN3(\FIFO[125][11] ), .IN4(n6732), 
        .Q(n542) );
  AO22X1 U5164 ( .IN1(n6960), .IN2(n6730), .IN3(\FIFO[125][12] ), .IN4(n6733), 
        .Q(n543) );
  AO22X1 U5165 ( .IN1(n6949), .IN2(n6730), .IN3(\FIFO[125][13] ), .IN4(n6733), 
        .Q(n544) );
  AO22X1 U5166 ( .IN1(n6938), .IN2(n6731), .IN3(\FIFO[125][14] ), .IN4(n6733), 
        .Q(n545) );
  AO22X1 U5167 ( .IN1(n6927), .IN2(n6730), .IN3(\FIFO[125][15] ), .IN4(n6733), 
        .Q(n546) );
  AO22X1 U5168 ( .IN1(n6916), .IN2(n6729), .IN3(\FIFO[125][16] ), .IN4(n6733), 
        .Q(n547) );
  AO22X1 U5169 ( .IN1(n6905), .IN2(n6731), .IN3(\FIFO[125][17] ), .IN4(n6733), 
        .Q(n548) );
  AO22X1 U5170 ( .IN1(n6894), .IN2(n6730), .IN3(\FIFO[125][18] ), .IN4(n6733), 
        .Q(n549) );
  AO22X1 U5171 ( .IN1(n6883), .IN2(n6729), .IN3(\FIFO[125][19] ), .IN4(n6733), 
        .Q(n550) );
  AO22X1 U5172 ( .IN1(n6872), .IN2(n6731), .IN3(\FIFO[125][20] ), .IN4(n6733), 
        .Q(n551) );
  AO22X1 U5173 ( .IN1(n6861), .IN2(n6729), .IN3(\FIFO[125][21] ), .IN4(n6733), 
        .Q(n552) );
  AO22X1 U5174 ( .IN1(n6850), .IN2(n6729), .IN3(\FIFO[125][22] ), .IN4(n6733), 
        .Q(n553) );
  AO22X1 U5175 ( .IN1(n6839), .IN2(n6729), .IN3(\FIFO[125][23] ), .IN4(n6733), 
        .Q(n554) );
  AO22X1 U5176 ( .IN1(n7098), .IN2(n6725), .IN3(\FIFO[124][0] ), .IN4(n6726), 
        .Q(n563) );
  AO22X1 U5177 ( .IN1(n7081), .IN2(n6725), .IN3(\FIFO[124][1] ), .IN4(n6726), 
        .Q(n564) );
  AO22X1 U5178 ( .IN1(n7070), .IN2(n6725), .IN3(\FIFO[124][2] ), .IN4(n6726), 
        .Q(n565) );
  AO22X1 U5179 ( .IN1(n7059), .IN2(n6725), .IN3(\FIFO[124][3] ), .IN4(n6726), 
        .Q(n566) );
  AO22X1 U5180 ( .IN1(n7048), .IN2(n6725), .IN3(\FIFO[124][4] ), .IN4(n6726), 
        .Q(n567) );
  AO22X1 U5181 ( .IN1(n7037), .IN2(n6725), .IN3(\FIFO[124][5] ), .IN4(n6726), 
        .Q(n568) );
  AO22X1 U5182 ( .IN1(n7026), .IN2(n6725), .IN3(\FIFO[124][6] ), .IN4(n6726), 
        .Q(n569) );
  AO22X1 U5183 ( .IN1(n7015), .IN2(n6724), .IN3(\FIFO[124][7] ), .IN4(n6726), 
        .Q(n570) );
  AO22X1 U5184 ( .IN1(n7004), .IN2(n6724), .IN3(\FIFO[124][8] ), .IN4(n6726), 
        .Q(n571) );
  AO22X1 U5185 ( .IN1(n6993), .IN2(n6724), .IN3(\FIFO[124][9] ), .IN4(n6726), 
        .Q(n572) );
  AO22X1 U5186 ( .IN1(n6982), .IN2(n6724), .IN3(\FIFO[124][10] ), .IN4(n6726), 
        .Q(n573) );
  AO22X1 U5187 ( .IN1(n6971), .IN2(n6724), .IN3(\FIFO[124][11] ), .IN4(n6726), 
        .Q(n574) );
  AO22X1 U5188 ( .IN1(n6894), .IN2(n6723), .IN3(\FIFO[124][18] ), .IN4(n6727), 
        .Q(n581) );
  AO22X1 U5189 ( .IN1(n6883), .IN2(n6723), .IN3(\FIFO[124][19] ), .IN4(n6727), 
        .Q(n582) );
  AO22X1 U5190 ( .IN1(n6872), .IN2(n6723), .IN3(\FIFO[124][20] ), .IN4(n6727), 
        .Q(n583) );
  AO22X1 U5191 ( .IN1(n6861), .IN2(n6725), .IN3(\FIFO[124][21] ), .IN4(n6727), 
        .Q(n584) );
  AO22X1 U5192 ( .IN1(n6850), .IN2(n6724), .IN3(\FIFO[124][22] ), .IN4(n6727), 
        .Q(n585) );
  AO22X1 U5193 ( .IN1(n6839), .IN2(n6723), .IN3(\FIFO[124][23] ), .IN4(n6727), 
        .Q(n586) );
  AO22X1 U5194 ( .IN1(n7098), .IN2(n6719), .IN3(\FIFO[123][0] ), .IN4(n6720), 
        .Q(n595) );
  AO22X1 U5195 ( .IN1(n7081), .IN2(n6719), .IN3(\FIFO[123][1] ), .IN4(n6720), 
        .Q(n596) );
  AO22X1 U5196 ( .IN1(n7070), .IN2(n6719), .IN3(\FIFO[123][2] ), .IN4(n6720), 
        .Q(n597) );
  AO22X1 U5197 ( .IN1(n7059), .IN2(n6719), .IN3(\FIFO[123][3] ), .IN4(n6720), 
        .Q(n598) );
  AO22X1 U5198 ( .IN1(n7048), .IN2(n6719), .IN3(\FIFO[123][4] ), .IN4(n6720), 
        .Q(n599) );
  AO22X1 U5199 ( .IN1(n7037), .IN2(n6719), .IN3(\FIFO[123][5] ), .IN4(n6720), 
        .Q(n600) );
  AO22X1 U5200 ( .IN1(n7026), .IN2(n6719), .IN3(\FIFO[123][6] ), .IN4(n6720), 
        .Q(n601) );
  AO22X1 U5201 ( .IN1(n7015), .IN2(n6718), .IN3(\FIFO[123][7] ), .IN4(n6720), 
        .Q(n602) );
  AO22X1 U5202 ( .IN1(n7004), .IN2(n6718), .IN3(\FIFO[123][8] ), .IN4(n6720), 
        .Q(n603) );
  AO22X1 U5203 ( .IN1(n6993), .IN2(n6718), .IN3(\FIFO[123][9] ), .IN4(n6720), 
        .Q(n604) );
  AO22X1 U5204 ( .IN1(n6982), .IN2(n6718), .IN3(\FIFO[123][10] ), .IN4(n6720), 
        .Q(n605) );
  AO22X1 U5205 ( .IN1(n6971), .IN2(n6718), .IN3(\FIFO[123][11] ), .IN4(n6720), 
        .Q(n606) );
  AO22X1 U5206 ( .IN1(n6960), .IN2(n6718), .IN3(\FIFO[123][12] ), .IN4(n6721), 
        .Q(n607) );
  AO22X1 U5207 ( .IN1(n6949), .IN2(n6718), .IN3(\FIFO[123][13] ), .IN4(n6721), 
        .Q(n608) );
  AO22X1 U5208 ( .IN1(n6938), .IN2(n6717), .IN3(\FIFO[123][14] ), .IN4(n6721), 
        .Q(n609) );
  AO22X1 U5209 ( .IN1(n6927), .IN2(n6717), .IN3(\FIFO[123][15] ), .IN4(n6721), 
        .Q(n610) );
  AO22X1 U5210 ( .IN1(n6916), .IN2(n6717), .IN3(\FIFO[123][16] ), .IN4(n6721), 
        .Q(n611) );
  AO22X1 U5211 ( .IN1(n6905), .IN2(n6717), .IN3(\FIFO[123][17] ), .IN4(n6721), 
        .Q(n612) );
  AO22X1 U5212 ( .IN1(n6894), .IN2(n6717), .IN3(\FIFO[123][18] ), .IN4(n6721), 
        .Q(n613) );
  AO22X1 U5213 ( .IN1(n6883), .IN2(n6717), .IN3(\FIFO[123][19] ), .IN4(n6721), 
        .Q(n614) );
  AO22X1 U5214 ( .IN1(n6872), .IN2(n6717), .IN3(\FIFO[123][20] ), .IN4(n6721), 
        .Q(n615) );
  AO22X1 U5215 ( .IN1(n6861), .IN2(n246), .IN3(\FIFO[123][21] ), .IN4(n6721), 
        .Q(n616) );
  AO22X1 U5216 ( .IN1(n6850), .IN2(n6719), .IN3(\FIFO[123][22] ), .IN4(n6721), 
        .Q(n617) );
  AO22X1 U5217 ( .IN1(n6839), .IN2(n6718), .IN3(\FIFO[123][23] ), .IN4(n6721), 
        .Q(n618) );
  AO22X1 U5218 ( .IN1(n7098), .IN2(n6713), .IN3(\FIFO[122][0] ), .IN4(n6714), 
        .Q(n627) );
  AO22X1 U5219 ( .IN1(n7081), .IN2(n6713), .IN3(\FIFO[122][1] ), .IN4(n6714), 
        .Q(n628) );
  AO22X1 U5220 ( .IN1(n7070), .IN2(n6713), .IN3(\FIFO[122][2] ), .IN4(n6714), 
        .Q(n629) );
  AO22X1 U5221 ( .IN1(n7059), .IN2(n6713), .IN3(\FIFO[122][3] ), .IN4(n6714), 
        .Q(n630) );
  AO22X1 U5222 ( .IN1(n7048), .IN2(n6713), .IN3(\FIFO[122][4] ), .IN4(n6714), 
        .Q(n631) );
  AO22X1 U5223 ( .IN1(n7037), .IN2(n6713), .IN3(\FIFO[122][5] ), .IN4(n6714), 
        .Q(n632) );
  AO22X1 U5224 ( .IN1(n7026), .IN2(n6713), .IN3(\FIFO[122][6] ), .IN4(n6714), 
        .Q(n633) );
  AO22X1 U5225 ( .IN1(n7015), .IN2(n6712), .IN3(\FIFO[122][7] ), .IN4(n6714), 
        .Q(n634) );
  AO22X1 U5226 ( .IN1(n7004), .IN2(n6712), .IN3(\FIFO[122][8] ), .IN4(n6714), 
        .Q(n635) );
  AO22X1 U5227 ( .IN1(n6993), .IN2(n6712), .IN3(\FIFO[122][9] ), .IN4(n6714), 
        .Q(n636) );
  AO22X1 U5228 ( .IN1(n6982), .IN2(n6712), .IN3(\FIFO[122][10] ), .IN4(n6714), 
        .Q(n637) );
  AO22X1 U5229 ( .IN1(n6971), .IN2(n6712), .IN3(\FIFO[122][11] ), .IN4(n6714), 
        .Q(n638) );
  AO22X1 U5230 ( .IN1(n6960), .IN2(n6712), .IN3(\FIFO[122][12] ), .IN4(n6715), 
        .Q(n639) );
  AO22X1 U5231 ( .IN1(n6949), .IN2(n6712), .IN3(\FIFO[122][13] ), .IN4(n6715), 
        .Q(n640) );
  AO22X1 U5232 ( .IN1(n6938), .IN2(n6711), .IN3(\FIFO[122][14] ), .IN4(n6715), 
        .Q(n641) );
  AO22X1 U5233 ( .IN1(n6927), .IN2(n6711), .IN3(\FIFO[122][15] ), .IN4(n6715), 
        .Q(n642) );
  AO22X1 U5234 ( .IN1(n6916), .IN2(n6711), .IN3(\FIFO[122][16] ), .IN4(n6715), 
        .Q(n643) );
  AO22X1 U5235 ( .IN1(n6905), .IN2(n6711), .IN3(\FIFO[122][17] ), .IN4(n6715), 
        .Q(n644) );
  AO22X1 U5236 ( .IN1(n6894), .IN2(n6711), .IN3(\FIFO[122][18] ), .IN4(n6715), 
        .Q(n645) );
  AO22X1 U5237 ( .IN1(n6883), .IN2(n6711), .IN3(\FIFO[122][19] ), .IN4(n6715), 
        .Q(n646) );
  AO22X1 U5238 ( .IN1(n6872), .IN2(n6711), .IN3(\FIFO[122][20] ), .IN4(n6715), 
        .Q(n647) );
  AO22X1 U5239 ( .IN1(n6861), .IN2(n6713), .IN3(\FIFO[122][21] ), .IN4(n6715), 
        .Q(n648) );
  AO22X1 U5240 ( .IN1(n6850), .IN2(n6712), .IN3(\FIFO[122][22] ), .IN4(n6715), 
        .Q(n649) );
  AO22X1 U5241 ( .IN1(n6839), .IN2(n6711), .IN3(\FIFO[122][23] ), .IN4(n6715), 
        .Q(n650) );
  AND2X1 U5242 ( .IN1(n53), .IN2(sync_flush), .Q(n204) );
  OR4X1 U5243 ( .IN1(n400), .IN2(n401), .IN3(N20), .IN4(N19), .Q(n53) );
  NBUFFX2 U5244 ( .INP(N15), .Z(n5972) );
  NBUFFX2 U5245 ( .INP(N15), .Z(n5971) );
  NBUFFX2 U5246 ( .INP(N15), .Z(n5970) );
  NBUFFX2 U5247 ( .INP(N15), .Z(n5969) );
  NBUFFX2 U5248 ( .INP(N15), .Z(n5968) );
  NBUFFX2 U5249 ( .INP(N15), .Z(n5967) );
  NBUFFX2 U5250 ( .INP(N15), .Z(n5966) );
  NBUFFX2 U5251 ( .INP(N15), .Z(n5965) );
  NBUFFX2 U5252 ( .INP(N16), .Z(n5788) );
  NBUFFX2 U5253 ( .INP(N16), .Z(n5787) );
  NBUFFX2 U5254 ( .INP(N16), .Z(n5786) );
  NBUFFX2 U5255 ( .INP(N16), .Z(n5785) );
  NBUFFX2 U5256 ( .INP(N16), .Z(n5784) );
  NBUFFX2 U5257 ( .INP(N16), .Z(n5783) );
  NBUFFX2 U5258 ( .INP(N16), .Z(n5782) );
  NBUFFX2 U5259 ( .INP(N17), .Z(n5776) );
  NBUFFX2 U5260 ( .INP(N17), .Z(n5777) );
  NBUFFX2 U5261 ( .INP(N17), .Z(n5778) );
  NBUFFX2 U5262 ( .INP(N17), .Z(n5779) );
  NBUFFX2 U5263 ( .INP(N17), .Z(n5780) );
  NBUFFX2 U5264 ( .INP(N17), .Z(n5781) );
  NBUFFX2 U5265 ( .INP(N18), .Z(n5756) );
  NBUFFX2 U5266 ( .INP(N18), .Z(n5757) );
  NBUFFX4 U5267 ( .INP(N19), .Z(n5730) );
  NBUFFX4 U5268 ( .INP(N19), .Z(n5731) );
  NBUFFX4 U5269 ( .INP(N19), .Z(n5732) );
  NBUFFX4 U5270 ( .INP(N19), .Z(n5733) );
  NBUFFX4 U5271 ( .INP(N19), .Z(n5734) );
  NBUFFX2 U5272 ( .INP(N20), .Z(n5726) );
  NBUFFX2 U5273 ( .INP(N20), .Z(n5727) );
  NBUFFX2 U5274 ( .INP(N20), .Z(n5728) );
  NBUFFX2 U5275 ( .INP(N20), .Z(n5729) );
  NBUFFX2 U5276 ( .INP(n5775), .Z(n5758) );
  NBUFFX2 U5277 ( .INP(N17), .Z(n5775) );
  NBUFFX2 U5278 ( .INP(N20), .Z(n5725) );
  NBUFFX2 U5279 ( .INP(N21), .Z(n5723) );
  NBUFFX2 U5280 ( .INP(N21), .Z(n5724) );
  NBUFFX4 U5281 ( .INP(flush), .Z(n7360) );
  NBUFFX4 U5282 ( .INP(flush), .Z(n7361) );
  NBUFFX2 U5283 ( .INP(flush), .Z(n7359) );
  OR2X1 U5284 ( .IN1(n7104), .IN2(\FIFO[0][0] ), .Q(n54) );
  OR2X1 U5285 ( .IN1(n7104), .IN2(\FIFO[0][1] ), .Q(n55) );
  OR2X1 U5286 ( .IN1(n7104), .IN2(\FIFO[0][2] ), .Q(n56) );
  OR2X1 U5287 ( .IN1(n7104), .IN2(\FIFO[0][3] ), .Q(n57) );
  OR2X1 U5288 ( .IN1(n7104), .IN2(\FIFO[0][4] ), .Q(n58) );
  OR2X1 U5289 ( .IN1(n7104), .IN2(\FIFO[0][5] ), .Q(n59) );
  OR2X1 U5290 ( .IN1(n7104), .IN2(\FIFO[0][6] ), .Q(n60) );
  OR2X1 U5291 ( .IN1(n7104), .IN2(\FIFO[0][7] ), .Q(n61) );
  OR2X1 U5292 ( .IN1(n7104), .IN2(\FIFO[0][8] ), .Q(n62) );
  OR2X1 U5293 ( .IN1(n7105), .IN2(\FIFO[0][12] ), .Q(n66) );
  OR2X1 U5294 ( .IN1(n7105), .IN2(\FIFO[0][13] ), .Q(n67) );
  OR2X1 U5295 ( .IN1(n7105), .IN2(\FIFO[0][14] ), .Q(n68) );
  OR2X1 U5296 ( .IN1(n7105), .IN2(\FIFO[0][15] ), .Q(n69) );
  OR2X1 U5297 ( .IN1(n7105), .IN2(\FIFO[0][16] ), .Q(n70) );
  OR2X1 U5298 ( .IN1(n7105), .IN2(\FIFO[0][17] ), .Q(n71) );
  OR2X1 U5299 ( .IN1(n7105), .IN2(\FIFO[0][18] ), .Q(n72) );
  OR2X1 U5300 ( .IN1(n7105), .IN2(\FIFO[0][19] ), .Q(n73) );
  OR2X1 U5301 ( .IN1(n7106), .IN2(\FIFO[0][24] ), .Q(n78) );
  OR2X1 U5302 ( .IN1(n7106), .IN2(\FIFO[0][25] ), .Q(n79) );
  OR2X1 U5303 ( .IN1(n7106), .IN2(\FIFO[0][26] ), .Q(n80) );
  OR2X1 U5304 ( .IN1(n7106), .IN2(\FIFO[0][28] ), .Q(n82) );
  NAND2X1 U5305 ( .IN1(n7354), .IN2(\FIFO[0][0] ), .QN(n86) );
  NAND2X1 U5306 ( .IN1(n7348), .IN2(\FIFO[0][1] ), .QN(n87) );
  NAND2X1 U5307 ( .IN1(n7341), .IN2(\FIFO[0][2] ), .QN(n88) );
  NAND2X1 U5308 ( .IN1(n7337), .IN2(\FIFO[0][6] ), .QN(n92) );
  NAND2X1 U5309 ( .IN1(n7357), .IN2(\FIFO[0][7] ), .QN(n93) );
  NAND2X1 U5310 ( .IN1(n7334), .IN2(\FIFO[0][8] ), .QN(n94) );
  NAND2X1 U5311 ( .IN1(n7351), .IN2(\FIFO[0][9] ), .QN(n95) );
  NAND2X1 U5312 ( .IN1(n7345), .IN2(\FIFO[0][10] ), .QN(n96) );
  NAND2X1 U5313 ( .IN1(n7358), .IN2(\FIFO[0][11] ), .QN(n97) );
  NAND2X1 U5314 ( .IN1(n7355), .IN2(\FIFO[0][12] ), .QN(n98) );
  NAND2X1 U5315 ( .IN1(n7357), .IN2(\FIFO[0][13] ), .QN(n99) );
  NAND2X1 U5316 ( .IN1(n7353), .IN2(\FIFO[0][14] ), .QN(n100) );
  NAND2X1 U5317 ( .IN1(n7358), .IN2(\FIFO[0][15] ), .QN(n101) );
  NAND2X1 U5318 ( .IN1(n7353), .IN2(\FIFO[0][16] ), .QN(n102) );
  NAND2X1 U5319 ( .IN1(n7334), .IN2(\FIFO[0][17] ), .QN(n103) );
  NAND2X1 U5320 ( .IN1(n7337), .IN2(\FIFO[0][20] ), .QN(n106) );
  NAND2X1 U5321 ( .IN1(n7348), .IN2(\FIFO[0][22] ), .QN(n108) );
  NAND2X1 U5322 ( .IN1(n7349), .IN2(\FIFO[0][23] ), .QN(n109) );
  NAND2X1 U5323 ( .IN1(n7350), .IN2(\FIFO[0][24] ), .QN(n110) );
  NAND2X1 U5324 ( .IN1(n7351), .IN2(\FIFO[0][25] ), .QN(n111) );
  NAND2X1 U5325 ( .IN1(n7344), .IN2(\FIFO[0][27] ), .QN(n113) );
  NAND2X1 U5326 ( .IN1(n7345), .IN2(\FIFO[0][29] ), .QN(n115) );
  NAND2X1 U5327 ( .IN1(n7346), .IN2(\FIFO[0][30] ), .QN(n116) );
  NAND2X1 U5328 ( .IN1(n7357), .IN2(\FIFO[0][31] ), .QN(n117) );
  MUX41X1 U5329 ( .IN1(\FIFO[124][0] ), .IN3(\FIFO[126][0] ), .IN2(
        \FIFO[125][0] ), .IN4(\FIFO[127][0] ), .S0(n5789), .S1(n5880), .Q(n118) );
  MUX41X1 U5330 ( .IN1(\FIFO[120][0] ), .IN3(\FIFO[122][0] ), .IN2(
        \FIFO[121][0] ), .IN4(\FIFO[123][0] ), .S0(n5789), .S1(n5891), .Q(n119) );
  MUX41X1 U5331 ( .IN1(\FIFO[116][0] ), .IN3(\FIFO[118][0] ), .IN2(
        \FIFO[117][0] ), .IN4(\FIFO[119][0] ), .S0(n5789), .S1(n5895), .Q(n120) );
  MUX41X1 U5332 ( .IN1(\FIFO[112][0] ), .IN3(\FIFO[114][0] ), .IN2(
        \FIFO[113][0] ), .IN4(\FIFO[115][0] ), .S0(n5789), .S1(n5874), .Q(n121) );
  MUX41X1 U5333 ( .IN1(n121), .IN3(n119), .IN2(n120), .IN4(n118), .S0(n5735), 
        .S1(n5758), .Q(n122) );
  MUX41X1 U5334 ( .IN1(\FIFO[108][0] ), .IN3(\FIFO[110][0] ), .IN2(
        \FIFO[109][0] ), .IN4(\FIFO[111][0] ), .S0(n5790), .S1(n5884), .Q(n123) );
  MUX41X1 U5335 ( .IN1(\FIFO[104][0] ), .IN3(\FIFO[106][0] ), .IN2(
        \FIFO[105][0] ), .IN4(\FIFO[107][0] ), .S0(n5790), .S1(n5885), .Q(n124) );
  MUX41X1 U5336 ( .IN1(\FIFO[100][0] ), .IN3(\FIFO[102][0] ), .IN2(
        \FIFO[101][0] ), .IN4(\FIFO[103][0] ), .S0(n5790), .S1(n5888), .Q(n125) );
  MUX41X1 U5337 ( .IN1(\FIFO[96][0] ), .IN3(\FIFO[98][0] ), .IN2(\FIFO[97][0] ), .IN4(\FIFO[99][0] ), .S0(n5790), .S1(n5889), .Q(n126) );
  MUX41X1 U5338 ( .IN1(n126), .IN3(n124), .IN2(n125), .IN4(n123), .S0(n5735), 
        .S1(n5758), .Q(n127) );
  MUX41X1 U5339 ( .IN1(\FIFO[92][0] ), .IN3(\FIFO[94][0] ), .IN2(\FIFO[93][0] ), .IN4(\FIFO[95][0] ), .S0(n5790), .S1(n5894), .Q(n128) );
  MUX41X1 U5340 ( .IN1(\FIFO[88][0] ), .IN3(\FIFO[90][0] ), .IN2(\FIFO[89][0] ), .IN4(\FIFO[91][0] ), .S0(n5790), .S1(n5887), .Q(n129) );
  MUX41X1 U5341 ( .IN1(\FIFO[84][0] ), .IN3(\FIFO[86][0] ), .IN2(\FIFO[85][0] ), .IN4(\FIFO[87][0] ), .S0(n5790), .S1(n5892), .Q(n130) );
  MUX41X1 U5342 ( .IN1(\FIFO[80][0] ), .IN3(\FIFO[82][0] ), .IN2(\FIFO[81][0] ), .IN4(\FIFO[83][0] ), .S0(n5790), .S1(n5893), .Q(n131) );
  MUX41X1 U5343 ( .IN1(n131), .IN3(n129), .IN2(n130), .IN4(n128), .S0(n5735), 
        .S1(n5758), .Q(n132) );
  MUX41X1 U5344 ( .IN1(\FIFO[76][0] ), .IN3(\FIFO[78][0] ), .IN2(\FIFO[77][0] ), .IN4(\FIFO[79][0] ), .S0(n5790), .S1(n5883), .Q(n133) );
  MUX41X1 U5345 ( .IN1(\FIFO[72][0] ), .IN3(\FIFO[74][0] ), .IN2(\FIFO[73][0] ), .IN4(\FIFO[75][0] ), .S0(n5790), .S1(n5896), .Q(n134) );
  MUX41X1 U5346 ( .IN1(\FIFO[68][0] ), .IN3(\FIFO[70][0] ), .IN2(\FIFO[69][0] ), .IN4(\FIFO[71][0] ), .S0(n5790), .S1(n5878), .Q(n135) );
  MUX41X1 U5347 ( .IN1(\FIFO[64][0] ), .IN3(\FIFO[66][0] ), .IN2(\FIFO[65][0] ), .IN4(\FIFO[67][0] ), .S0(n5790), .S1(n5881), .Q(n136) );
  MUX41X1 U5348 ( .IN1(n136), .IN3(n134), .IN2(n135), .IN4(n133), .S0(n5735), 
        .S1(n5758), .Q(n137) );
  MUX41X1 U5349 ( .IN1(n137), .IN3(n127), .IN2(n132), .IN4(n122), .S0(n5725), 
        .S1(N19), .Q(n138) );
  MUX41X1 U5350 ( .IN1(\FIFO[60][0] ), .IN3(\FIFO[62][0] ), .IN2(\FIFO[61][0] ), .IN4(\FIFO[63][0] ), .S0(n5791), .S1(n5883), .Q(n139) );
  MUX41X1 U5351 ( .IN1(\FIFO[56][0] ), .IN3(\FIFO[58][0] ), .IN2(\FIFO[57][0] ), .IN4(\FIFO[59][0] ), .S0(n5791), .S1(n5888), .Q(n140) );
  MUX41X1 U5352 ( .IN1(\FIFO[52][0] ), .IN3(\FIFO[54][0] ), .IN2(\FIFO[53][0] ), .IN4(\FIFO[55][0] ), .S0(n5791), .S1(n5878), .Q(n141) );
  MUX41X1 U5353 ( .IN1(\FIFO[48][0] ), .IN3(\FIFO[50][0] ), .IN2(\FIFO[49][0] ), .IN4(\FIFO[51][0] ), .S0(n5791), .S1(n5881), .Q(n142) );
  MUX41X1 U5354 ( .IN1(n142), .IN3(n140), .IN2(n141), .IN4(n139), .S0(n5736), 
        .S1(n5779), .Q(n143) );
  MUX41X1 U5355 ( .IN1(\FIFO[44][0] ), .IN3(\FIFO[46][0] ), .IN2(\FIFO[45][0] ), .IN4(\FIFO[47][0] ), .S0(n5791), .S1(n5887), .Q(n144) );
  MUX41X1 U5356 ( .IN1(\FIFO[40][0] ), .IN3(\FIFO[42][0] ), .IN2(\FIFO[41][0] ), .IN4(\FIFO[43][0] ), .S0(n5791), .S1(n5889), .Q(n145) );
  MUX41X1 U5357 ( .IN1(\FIFO[36][0] ), .IN3(\FIFO[38][0] ), .IN2(\FIFO[37][0] ), .IN4(\FIFO[39][0] ), .S0(n5791), .S1(n5885), .Q(n146) );
  MUX41X1 U5358 ( .IN1(\FIFO[32][0] ), .IN3(\FIFO[34][0] ), .IN2(\FIFO[33][0] ), .IN4(\FIFO[35][0] ), .S0(n5791), .S1(n5886), .Q(n147) );
  MUX41X1 U5359 ( .IN1(n147), .IN3(n145), .IN2(n146), .IN4(n144), .S0(n5736), 
        .S1(n5780), .Q(n148) );
  MUX41X1 U5360 ( .IN1(\FIFO[28][0] ), .IN3(\FIFO[30][0] ), .IN2(\FIFO[29][0] ), .IN4(\FIFO[31][0] ), .S0(n5791), .S1(n5894), .Q(n149) );
  MUX41X1 U5361 ( .IN1(\FIFO[24][0] ), .IN3(\FIFO[26][0] ), .IN2(\FIFO[25][0] ), .IN4(\FIFO[27][0] ), .S0(n5791), .S1(n5884), .Q(n150) );
  MUX41X1 U5362 ( .IN1(\FIFO[20][0] ), .IN3(\FIFO[22][0] ), .IN2(\FIFO[21][0] ), .IN4(\FIFO[23][0] ), .S0(n5791), .S1(n5892), .Q(n151) );
  MUX41X1 U5363 ( .IN1(\FIFO[16][0] ), .IN3(\FIFO[18][0] ), .IN2(\FIFO[17][0] ), .IN4(\FIFO[19][0] ), .S0(n5791), .S1(n5893), .Q(n152) );
  MUX41X1 U5364 ( .IN1(n152), .IN3(n150), .IN2(n151), .IN4(n149), .S0(n5736), 
        .S1(n5781), .Q(n153) );
  MUX41X1 U5365 ( .IN1(\FIFO[12][0] ), .IN3(\FIFO[14][0] ), .IN2(\FIFO[13][0] ), .IN4(\FIFO[15][0] ), .S0(n5792), .S1(n5893), .Q(n154) );
  MUX41X1 U5366 ( .IN1(\FIFO[8][0] ), .IN3(\FIFO[10][0] ), .IN2(\FIFO[9][0] ), 
        .IN4(\FIFO[11][0] ), .S0(n5792), .S1(n5878), .Q(n155) );
  MUX41X1 U5367 ( .IN1(\FIFO[4][0] ), .IN3(\FIFO[6][0] ), .IN2(\FIFO[5][0] ), 
        .IN4(\FIFO[7][0] ), .S0(n5792), .S1(n5891), .Q(n156) );
  MUX41X1 U5368 ( .IN1(\FIFO[0][0] ), .IN3(\FIFO[2][0] ), .IN2(\FIFO[1][0] ), 
        .IN4(\FIFO[3][0] ), .S0(n5792), .S1(n5892), .Q(n157) );
  MUX41X1 U5369 ( .IN1(n157), .IN3(n155), .IN2(n156), .IN4(n154), .S0(n5736), 
        .S1(n5777), .Q(n158) );
  MUX41X1 U5370 ( .IN1(n158), .IN3(n148), .IN2(n153), .IN4(n143), .S0(n5725), 
        .S1(N19), .Q(n159) );
  MUX21X1 U5371 ( .IN1(n159), .IN2(n138), .S(N21), .Q(N250) );
  MUX41X1 U5372 ( .IN1(\FIFO[124][1] ), .IN3(\FIFO[126][1] ), .IN2(
        \FIFO[125][1] ), .IN4(\FIFO[127][1] ), .S0(n5792), .S1(n5883), .Q(n160) );
  MUX41X1 U5373 ( .IN1(\FIFO[120][1] ), .IN3(\FIFO[122][1] ), .IN2(
        \FIFO[121][1] ), .IN4(\FIFO[123][1] ), .S0(n5792), .S1(n5887), .Q(n161) );
  MUX41X1 U5374 ( .IN1(\FIFO[116][1] ), .IN3(\FIFO[118][1] ), .IN2(
        \FIFO[117][1] ), .IN4(\FIFO[119][1] ), .S0(n5792), .S1(n5894), .Q(n162) );
  MUX41X1 U5375 ( .IN1(\FIFO[112][1] ), .IN3(\FIFO[114][1] ), .IN2(
        \FIFO[113][1] ), .IN4(\FIFO[115][1] ), .S0(n5792), .S1(n5881), .Q(n163) );
  MUX41X1 U5376 ( .IN1(n163), .IN3(n161), .IN2(n162), .IN4(n160), .S0(n5736), 
        .S1(n5778), .Q(n164) );
  MUX41X1 U5377 ( .IN1(\FIFO[108][1] ), .IN3(\FIFO[110][1] ), .IN2(
        \FIFO[109][1] ), .IN4(\FIFO[111][1] ), .S0(n5792), .S1(n5886), .Q(n165) );
  MUX41X1 U5378 ( .IN1(\FIFO[104][1] ), .IN3(\FIFO[106][1] ), .IN2(
        \FIFO[105][1] ), .IN4(\FIFO[107][1] ), .S0(n5792), .S1(n5965), .Q(n166) );
  MUX41X1 U5379 ( .IN1(\FIFO[100][1] ), .IN3(\FIFO[102][1] ), .IN2(
        \FIFO[101][1] ), .IN4(\FIFO[103][1] ), .S0(n5792), .S1(n5884), .Q(n167) );
  MUX41X1 U5380 ( .IN1(\FIFO[96][1] ), .IN3(\FIFO[98][1] ), .IN2(\FIFO[97][1] ), .IN4(\FIFO[99][1] ), .S0(n5792), .S1(n5885), .Q(n168) );
  MUX41X1 U5381 ( .IN1(n168), .IN3(n166), .IN2(n167), .IN4(n165), .S0(n5736), 
        .S1(n5779), .Q(n169) );
  MUX41X1 U5382 ( .IN1(\FIFO[92][1] ), .IN3(\FIFO[94][1] ), .IN2(\FIFO[93][1] ), .IN4(\FIFO[95][1] ), .S0(n5793), .S1(n5876), .Q(n170) );
  MUX41X1 U5383 ( .IN1(\FIFO[88][1] ), .IN3(\FIFO[90][1] ), .IN2(\FIFO[89][1] ), .IN4(\FIFO[91][1] ), .S0(n5793), .S1(n5879), .Q(n171) );
  MUX41X1 U5384 ( .IN1(\FIFO[84][1] ), .IN3(\FIFO[86][1] ), .IN2(\FIFO[85][1] ), .IN4(\FIFO[87][1] ), .S0(n5793), .S1(n5892), .Q(n172) );
  MUX41X1 U5385 ( .IN1(\FIFO[80][1] ), .IN3(\FIFO[82][1] ), .IN2(\FIFO[81][1] ), .IN4(\FIFO[83][1] ), .S0(n5793), .S1(n5896), .Q(n173) );
  MUX41X1 U5386 ( .IN1(n173), .IN3(n171), .IN2(n172), .IN4(n170), .S0(n5736), 
        .S1(n5776), .Q(n174) );
  MUX41X1 U5387 ( .IN1(\FIFO[76][1] ), .IN3(\FIFO[78][1] ), .IN2(\FIFO[77][1] ), .IN4(\FIFO[79][1] ), .S0(n5793), .S1(n5874), .Q(n175) );
  MUX41X1 U5388 ( .IN1(\FIFO[72][1] ), .IN3(\FIFO[74][1] ), .IN2(\FIFO[73][1] ), .IN4(\FIFO[75][1] ), .S0(n5793), .S1(n5890), .Q(n176) );
  MUX41X1 U5389 ( .IN1(\FIFO[68][1] ), .IN3(\FIFO[70][1] ), .IN2(\FIFO[69][1] ), .IN4(\FIFO[71][1] ), .S0(n5793), .S1(n5965), .Q(n177) );
  MUX41X1 U5390 ( .IN1(\FIFO[64][1] ), .IN3(\FIFO[66][1] ), .IN2(\FIFO[65][1] ), .IN4(\FIFO[67][1] ), .S0(n5793), .S1(n5882), .Q(n178) );
  MUX41X1 U5391 ( .IN1(n178), .IN3(n176), .IN2(n177), .IN4(n175), .S0(n5736), 
        .S1(n5777), .Q(n179) );
  MUX41X1 U5392 ( .IN1(n179), .IN3(n169), .IN2(n174), .IN4(n164), .S0(n5725), 
        .S1(N19), .Q(n180) );
  MUX41X1 U5393 ( .IN1(\FIFO[60][1] ), .IN3(\FIFO[62][1] ), .IN2(\FIFO[61][1] ), .IN4(\FIFO[63][1] ), .S0(n5793), .S1(n5876), .Q(n181) );
  MUX41X1 U5394 ( .IN1(\FIFO[56][1] ), .IN3(\FIFO[58][1] ), .IN2(\FIFO[57][1] ), .IN4(\FIFO[59][1] ), .S0(n5793), .S1(n5880), .Q(n182) );
  MUX41X1 U5395 ( .IN1(\FIFO[52][1] ), .IN3(\FIFO[54][1] ), .IN2(\FIFO[53][1] ), .IN4(\FIFO[55][1] ), .S0(n5793), .S1(n5971), .Q(n183) );
  MUX41X1 U5396 ( .IN1(\FIFO[48][1] ), .IN3(\FIFO[50][1] ), .IN2(\FIFO[49][1] ), .IN4(\FIFO[51][1] ), .S0(n5793), .S1(n5966), .Q(n184) );
  MUX41X1 U5397 ( .IN1(n184), .IN3(n182), .IN2(n183), .IN4(n181), .S0(n5736), 
        .S1(n5778), .Q(n185) );
  MUX41X1 U5398 ( .IN1(\FIFO[44][1] ), .IN3(\FIFO[46][1] ), .IN2(\FIFO[45][1] ), .IN4(\FIFO[47][1] ), .S0(n5789), .S1(n5888), .Q(n186) );
  MUX41X1 U5399 ( .IN1(\FIFO[40][1] ), .IN3(\FIFO[42][1] ), .IN2(\FIFO[41][1] ), .IN4(\FIFO[43][1] ), .S0(n5789), .S1(n5968), .Q(n187) );
  MUX41X1 U5400 ( .IN1(\FIFO[36][1] ), .IN3(\FIFO[38][1] ), .IN2(\FIFO[37][1] ), .IN4(\FIFO[39][1] ), .S0(n5789), .S1(n5885), .Q(n188) );
  MUX41X1 U5401 ( .IN1(\FIFO[32][1] ), .IN3(\FIFO[34][1] ), .IN2(\FIFO[33][1] ), .IN4(\FIFO[35][1] ), .S0(n5789), .S1(n5886), .Q(n189) );
  MUX41X1 U5402 ( .IN1(n189), .IN3(n187), .IN2(n188), .IN4(n186), .S0(n5736), 
        .S1(n5781), .Q(n190) );
  MUX41X1 U5403 ( .IN1(\FIFO[28][1] ), .IN3(\FIFO[30][1] ), .IN2(\FIFO[29][1] ), .IN4(\FIFO[31][1] ), .S0(n5841), .S1(n5889), .Q(n191) );
  MUX41X1 U5404 ( .IN1(\FIFO[24][1] ), .IN3(\FIFO[26][1] ), .IN2(\FIFO[25][1] ), .IN4(\FIFO[27][1] ), .S0(n5870), .S1(n5884), .Q(n192) );
  MUX41X1 U5405 ( .IN1(\FIFO[20][1] ), .IN3(\FIFO[22][1] ), .IN2(\FIFO[21][1] ), .IN4(\FIFO[23][1] ), .S0(n5814), .S1(n5893), .Q(n193) );
  MUX41X1 U5406 ( .IN1(\FIFO[16][1] ), .IN3(\FIFO[18][1] ), .IN2(\FIFO[17][1] ), .IN4(\FIFO[19][1] ), .S0(n5789), .S1(n5894), .Q(n194) );
  MUX41X1 U5407 ( .IN1(n194), .IN3(n192), .IN2(n193), .IN4(n191), .S0(n5736), 
        .S1(n5776), .Q(n195) );
  MUX41X1 U5408 ( .IN1(\FIFO[12][1] ), .IN3(\FIFO[14][1] ), .IN2(\FIFO[13][1] ), .IN4(\FIFO[15][1] ), .S0(n5789), .S1(n5883), .Q(n196) );
  MUX41X1 U5409 ( .IN1(\FIFO[8][1] ), .IN3(\FIFO[10][1] ), .IN2(\FIFO[9][1] ), 
        .IN4(\FIFO[11][1] ), .S0(n5789), .S1(n5887), .Q(n197) );
  MUX41X1 U5410 ( .IN1(\FIFO[4][1] ), .IN3(\FIFO[6][1] ), .IN2(\FIFO[5][1] ), 
        .IN4(\FIFO[7][1] ), .S0(n5789), .S1(n5878), .Q(n198) );
  MUX41X1 U5411 ( .IN1(\FIFO[0][1] ), .IN3(\FIFO[2][1] ), .IN2(\FIFO[1][1] ), 
        .IN4(\FIFO[3][1] ), .S0(n5838), .S1(n5881), .Q(n199) );
  MUX41X1 U5412 ( .IN1(n199), .IN3(n197), .IN2(n198), .IN4(n196), .S0(n5736), 
        .S1(n5780), .Q(n200) );
  MUX41X1 U5413 ( .IN1(n200), .IN3(n190), .IN2(n195), .IN4(n185), .S0(n5725), 
        .S1(N19), .Q(n201) );
  MUX21X1 U5414 ( .IN1(n201), .IN2(n180), .S(N21), .Q(N249) );
  MUX41X1 U5415 ( .IN1(\FIFO[124][2] ), .IN3(\FIFO[126][2] ), .IN2(
        \FIFO[125][2] ), .IN4(\FIFO[127][2] ), .S0(n5794), .S1(n5889), .Q(n202) );
  MUX41X1 U5416 ( .IN1(\FIFO[120][2] ), .IN3(\FIFO[122][2] ), .IN2(
        \FIFO[121][2] ), .IN4(\FIFO[123][2] ), .S0(n5794), .S1(n5890), .Q(n203) );
  MUX41X1 U5417 ( .IN1(\FIFO[116][2] ), .IN3(\FIFO[118][2] ), .IN2(
        \FIFO[117][2] ), .IN4(\FIFO[119][2] ), .S0(n5794), .S1(n5887), .Q(n205) );
  MUX41X1 U5418 ( .IN1(\FIFO[112][2] ), .IN3(\FIFO[114][2] ), .IN2(
        \FIFO[113][2] ), .IN4(\FIFO[115][2] ), .S0(n5794), .S1(n5888), .Q(n207) );
  MUX41X1 U5419 ( .IN1(n207), .IN3(n203), .IN2(n205), .IN4(n202), .S0(n5735), 
        .S1(n5778), .Q(n208) );
  MUX41X1 U5420 ( .IN1(\FIFO[108][2] ), .IN3(\FIFO[110][2] ), .IN2(
        \FIFO[109][2] ), .IN4(\FIFO[111][2] ), .S0(n5794), .S1(n5879), .Q(n209) );
  MUX41X1 U5421 ( .IN1(\FIFO[104][2] ), .IN3(\FIFO[106][2] ), .IN2(
        \FIFO[105][2] ), .IN4(\FIFO[107][2] ), .S0(n5794), .S1(n5877), .Q(n210) );
  MUX41X1 U5422 ( .IN1(\FIFO[100][2] ), .IN3(\FIFO[102][2] ), .IN2(
        \FIFO[101][2] ), .IN4(\FIFO[103][2] ), .S0(n5794), .S1(n5875), .Q(n211) );
  MUX41X1 U5423 ( .IN1(\FIFO[96][2] ), .IN3(\FIFO[98][2] ), .IN2(\FIFO[97][2] ), .IN4(\FIFO[99][2] ), .S0(n5794), .S1(n5882), .Q(n212) );
  MUX41X1 U5424 ( .IN1(n212), .IN3(n210), .IN2(n211), .IN4(n209), .S0(n5735), 
        .S1(n5776), .Q(n213) );
  MUX41X1 U5425 ( .IN1(\FIFO[92][2] ), .IN3(\FIFO[94][2] ), .IN2(\FIFO[93][2] ), .IN4(\FIFO[95][2] ), .S0(n5794), .S1(n5886), .Q(n214) );
  MUX41X1 U5426 ( .IN1(\FIFO[88][2] ), .IN3(\FIFO[90][2] ), .IN2(\FIFO[89][2] ), .IN4(\FIFO[91][2] ), .S0(n5794), .S1(n5967), .Q(n215) );
  MUX41X1 U5427 ( .IN1(\FIFO[84][2] ), .IN3(\FIFO[86][2] ), .IN2(\FIFO[85][2] ), .IN4(\FIFO[87][2] ), .S0(n5794), .S1(n5884), .Q(n216) );
  MUX41X1 U5428 ( .IN1(\FIFO[80][2] ), .IN3(\FIFO[82][2] ), .IN2(\FIFO[81][2] ), .IN4(\FIFO[83][2] ), .S0(n5794), .S1(n5885), .Q(n217) );
  MUX41X1 U5429 ( .IN1(n217), .IN3(n215), .IN2(n216), .IN4(n214), .S0(n5735), 
        .S1(N17), .Q(n218) );
  MUX41X1 U5430 ( .IN1(\FIFO[76][2] ), .IN3(\FIFO[78][2] ), .IN2(\FIFO[77][2] ), .IN4(\FIFO[79][2] ), .S0(n5795), .S1(n5881), .Q(n219) );
  MUX41X1 U5431 ( .IN1(\FIFO[72][2] ), .IN3(\FIFO[74][2] ), .IN2(\FIFO[73][2] ), .IN4(\FIFO[75][2] ), .S0(n5795), .S1(n5965), .Q(n220) );
  MUX41X1 U5432 ( .IN1(\FIFO[68][2] ), .IN3(\FIFO[70][2] ), .IN2(\FIFO[69][2] ), .IN4(\FIFO[71][2] ), .S0(n5795), .S1(n5891), .Q(n221) );
  MUX41X1 U5433 ( .IN1(\FIFO[64][2] ), .IN3(\FIFO[66][2] ), .IN2(\FIFO[65][2] ), .IN4(\FIFO[67][2] ), .S0(n5795), .S1(n5878), .Q(n222) );
  MUX41X1 U5434 ( .IN1(n222), .IN3(n220), .IN2(n221), .IN4(n219), .S0(n5735), 
        .S1(n5780), .Q(n223) );
  MUX41X1 U5435 ( .IN1(n223), .IN3(n213), .IN2(n218), .IN4(n208), .S0(n5726), 
        .S1(n5730), .Q(n224) );
  MUX41X1 U5436 ( .IN1(\FIFO[60][2] ), .IN3(\FIFO[62][2] ), .IN2(\FIFO[61][2] ), .IN4(\FIFO[63][2] ), .S0(n5795), .S1(n5879), .Q(n225) );
  MUX41X1 U5437 ( .IN1(\FIFO[56][2] ), .IN3(\FIFO[58][2] ), .IN2(\FIFO[57][2] ), .IN4(\FIFO[59][2] ), .S0(n5795), .S1(n5894), .Q(n226) );
  MUX41X1 U5438 ( .IN1(\FIFO[52][2] ), .IN3(\FIFO[54][2] ), .IN2(\FIFO[53][2] ), .IN4(\FIFO[55][2] ), .S0(n5795), .S1(n5880), .Q(n227) );
  MUX41X1 U5439 ( .IN1(\FIFO[48][2] ), .IN3(\FIFO[50][2] ), .IN2(\FIFO[49][2] ), .IN4(\FIFO[51][2] ), .S0(n5795), .S1(n5882), .Q(n228) );
  MUX41X1 U5440 ( .IN1(n228), .IN3(n226), .IN2(n227), .IN4(n225), .S0(n5756), 
        .S1(N17), .Q(n229) );
  MUX41X1 U5441 ( .IN1(\FIFO[44][2] ), .IN3(\FIFO[46][2] ), .IN2(\FIFO[45][2] ), .IN4(\FIFO[47][2] ), .S0(n5795), .S1(n5893), .Q(n230) );
  MUX41X1 U5442 ( .IN1(\FIFO[40][2] ), .IN3(\FIFO[42][2] ), .IN2(\FIFO[41][2] ), .IN4(\FIFO[43][2] ), .S0(n5795), .S1(n5883), .Q(n231) );
  MUX41X1 U5443 ( .IN1(\FIFO[36][2] ), .IN3(\FIFO[38][2] ), .IN2(\FIFO[37][2] ), .IN4(\FIFO[39][2] ), .S0(n5795), .S1(n5890), .Q(n232) );
  MUX41X1 U5444 ( .IN1(\FIFO[32][2] ), .IN3(\FIFO[34][2] ), .IN2(\FIFO[33][2] ), .IN4(\FIFO[35][2] ), .S0(n5795), .S1(n5892), .Q(n233) );
  MUX41X1 U5445 ( .IN1(n233), .IN3(n231), .IN2(n232), .IN4(n230), .S0(n5735), 
        .S1(n5776), .Q(n234) );
  MUX41X1 U5446 ( .IN1(\FIFO[28][2] ), .IN3(\FIFO[30][2] ), .IN2(\FIFO[29][2] ), .IN4(\FIFO[31][2] ), .S0(n5796), .S1(n5895), .Q(n235) );
  MUX41X1 U5447 ( .IN1(\FIFO[24][2] ), .IN3(\FIFO[26][2] ), .IN2(\FIFO[25][2] ), .IN4(\FIFO[27][2] ), .S0(n5796), .S1(n5966), .Q(n236) );
  MUX41X1 U5448 ( .IN1(\FIFO[20][2] ), .IN3(\FIFO[22][2] ), .IN2(\FIFO[21][2] ), .IN4(\FIFO[23][2] ), .S0(n5796), .S1(n5888), .Q(n237) );
  MUX41X1 U5449 ( .IN1(\FIFO[16][2] ), .IN3(\FIFO[18][2] ), .IN2(\FIFO[17][2] ), .IN4(\FIFO[19][2] ), .S0(n5796), .S1(n5889), .Q(n398) );
  MUX41X1 U5450 ( .IN1(n398), .IN3(n236), .IN2(n237), .IN4(n235), .S0(n5741), 
        .S1(n5779), .Q(n399) );
  MUX41X1 U5451 ( .IN1(\FIFO[12][2] ), .IN3(\FIFO[14][2] ), .IN2(\FIFO[13][2] ), .IN4(\FIFO[15][2] ), .S0(n5796), .S1(n5896), .Q(n402) );
  MUX41X1 U5452 ( .IN1(\FIFO[8][2] ), .IN3(\FIFO[10][2] ), .IN2(\FIFO[9][2] ), 
        .IN4(\FIFO[11][2] ), .S0(n5796), .S1(n5875), .Q(n403) );
  MUX41X1 U5453 ( .IN1(\FIFO[4][2] ), .IN3(\FIFO[6][2] ), .IN2(\FIFO[5][2] ), 
        .IN4(\FIFO[7][2] ), .S0(n5796), .S1(n5968), .Q(n404) );
  MUX41X1 U5454 ( .IN1(\FIFO[0][2] ), .IN3(\FIFO[2][2] ), .IN2(\FIFO[1][2] ), 
        .IN4(\FIFO[3][2] ), .S0(n5796), .S1(n5874), .Q(n405) );
  MUX41X1 U5455 ( .IN1(n405), .IN3(n403), .IN2(n404), .IN4(n402), .S0(n5740), 
        .S1(N17), .Q(n406) );
  MUX41X1 U5456 ( .IN1(n406), .IN3(n234), .IN2(n399), .IN4(n229), .S0(n5726), 
        .S1(n5730), .Q(n407) );
  MUX21X1 U5457 ( .IN1(n407), .IN2(n224), .S(N21), .Q(N248) );
  MUX41X1 U5458 ( .IN1(\FIFO[124][3] ), .IN3(\FIFO[126][3] ), .IN2(
        \FIFO[125][3] ), .IN4(\FIFO[127][3] ), .S0(n5796), .S1(n5877), .Q(n408) );
  MUX41X1 U5459 ( .IN1(\FIFO[120][3] ), .IN3(\FIFO[122][3] ), .IN2(
        \FIFO[121][3] ), .IN4(\FIFO[123][3] ), .S0(n5796), .S1(n5874), .Q(n409) );
  MUX41X1 U5460 ( .IN1(\FIFO[116][3] ), .IN3(\FIFO[118][3] ), .IN2(
        \FIFO[117][3] ), .IN4(\FIFO[119][3] ), .S0(n5796), .S1(n5895), .Q(n410) );
  MUX41X1 U5461 ( .IN1(\FIFO[112][3] ), .IN3(\FIFO[114][3] ), .IN2(
        \FIFO[113][3] ), .IN4(\FIFO[115][3] ), .S0(n5796), .S1(n5876), .Q(n411) );
  MUX41X1 U5462 ( .IN1(n411), .IN3(n409), .IN2(n410), .IN4(n408), .S0(n5735), 
        .S1(n5777), .Q(n412) );
  MUX41X1 U5463 ( .IN1(\FIFO[108][3] ), .IN3(\FIFO[110][3] ), .IN2(
        \FIFO[109][3] ), .IN4(\FIFO[111][3] ), .S0(n5797), .S1(n5892), .Q(n413) );
  MUX41X1 U5464 ( .IN1(\FIFO[104][3] ), .IN3(\FIFO[106][3] ), .IN2(
        \FIFO[105][3] ), .IN4(\FIFO[107][3] ), .S0(n5797), .S1(n5891), .Q(n414) );
  MUX41X1 U5465 ( .IN1(\FIFO[100][3] ), .IN3(\FIFO[102][3] ), .IN2(
        \FIFO[101][3] ), .IN4(\FIFO[103][3] ), .S0(n5797), .S1(n5879), .Q(n415) );
  MUX41X1 U5466 ( .IN1(\FIFO[96][3] ), .IN3(\FIFO[98][3] ), .IN2(\FIFO[97][3] ), .IN4(\FIFO[99][3] ), .S0(n5797), .S1(n5890), .Q(n416) );
  MUX41X1 U5467 ( .IN1(n416), .IN3(n414), .IN2(n415), .IN4(n413), .S0(n5735), 
        .S1(n5779), .Q(n417) );
  MUX41X1 U5468 ( .IN1(\FIFO[92][3] ), .IN3(\FIFO[94][3] ), .IN2(\FIFO[93][3] ), .IN4(\FIFO[95][3] ), .S0(n5797), .S1(n5877), .Q(n418) );
  MUX41X1 U5469 ( .IN1(\FIFO[88][3] ), .IN3(\FIFO[90][3] ), .IN2(\FIFO[89][3] ), .IN4(\FIFO[91][3] ), .S0(n5797), .S1(n5882), .Q(n419) );
  MUX41X1 U5470 ( .IN1(\FIFO[84][3] ), .IN3(\FIFO[86][3] ), .IN2(\FIFO[85][3] ), .IN4(\FIFO[87][3] ), .S0(n5797), .S1(n5877), .Q(n420) );
  MUX41X1 U5471 ( .IN1(\FIFO[80][3] ), .IN3(\FIFO[82][3] ), .IN2(\FIFO[81][3] ), .IN4(\FIFO[83][3] ), .S0(n5797), .S1(n5971), .Q(n421) );
  MUX41X1 U5472 ( .IN1(n421), .IN3(n419), .IN2(n420), .IN4(n418), .S0(n5756), 
        .S1(N17), .Q(n422) );
  MUX41X1 U5473 ( .IN1(\FIFO[76][3] ), .IN3(\FIFO[78][3] ), .IN2(\FIFO[77][3] ), .IN4(\FIFO[79][3] ), .S0(n5797), .S1(n5880), .Q(n423) );
  MUX41X1 U5474 ( .IN1(\FIFO[72][3] ), .IN3(\FIFO[74][3] ), .IN2(\FIFO[73][3] ), .IN4(\FIFO[75][3] ), .S0(n5797), .S1(n5891), .Q(n424) );
  MUX41X1 U5475 ( .IN1(\FIFO[68][3] ), .IN3(\FIFO[70][3] ), .IN2(\FIFO[69][3] ), .IN4(\FIFO[71][3] ), .S0(n5797), .S1(n5896), .Q(n425) );
  MUX41X1 U5476 ( .IN1(\FIFO[64][3] ), .IN3(\FIFO[66][3] ), .IN2(\FIFO[65][3] ), .IN4(\FIFO[67][3] ), .S0(n5797), .S1(n5895), .Q(n426) );
  MUX41X1 U5477 ( .IN1(n426), .IN3(n424), .IN2(n425), .IN4(n423), .S0(n5735), 
        .S1(n5781), .Q(n427) );
  MUX41X1 U5478 ( .IN1(n427), .IN3(n417), .IN2(n422), .IN4(n412), .S0(n5726), 
        .S1(n5730), .Q(n428) );
  MUX41X1 U5479 ( .IN1(\FIFO[60][3] ), .IN3(\FIFO[62][3] ), .IN2(\FIFO[61][3] ), .IN4(\FIFO[63][3] ), .S0(n5798), .S1(n5889), .Q(n429) );
  MUX41X1 U5480 ( .IN1(\FIFO[56][3] ), .IN3(\FIFO[58][3] ), .IN2(\FIFO[57][3] ), .IN4(\FIFO[59][3] ), .S0(n5798), .S1(n5875), .Q(n430) );
  MUX41X1 U5481 ( .IN1(\FIFO[52][3] ), .IN3(\FIFO[54][3] ), .IN2(\FIFO[53][3] ), .IN4(\FIFO[55][3] ), .S0(n5798), .S1(n5887), .Q(n431) );
  MUX41X1 U5482 ( .IN1(\FIFO[48][3] ), .IN3(\FIFO[50][3] ), .IN2(\FIFO[49][3] ), .IN4(\FIFO[51][3] ), .S0(n5798), .S1(n5888), .Q(n432) );
  MUX41X1 U5483 ( .IN1(n432), .IN3(n430), .IN2(n431), .IN4(n429), .S0(n5737), 
        .S1(n5778), .Q(n433) );
  MUX41X1 U5484 ( .IN1(\FIFO[44][3] ), .IN3(\FIFO[46][3] ), .IN2(\FIFO[45][3] ), .IN4(\FIFO[47][3] ), .S0(n5798), .S1(n5896), .Q(n434) );
  MUX41X1 U5485 ( .IN1(\FIFO[40][3] ), .IN3(\FIFO[42][3] ), .IN2(\FIFO[41][3] ), .IN4(\FIFO[43][3] ), .S0(n5798), .S1(n5876), .Q(n435) );
  MUX41X1 U5486 ( .IN1(\FIFO[36][3] ), .IN3(\FIFO[38][3] ), .IN2(\FIFO[37][3] ), .IN4(\FIFO[39][3] ), .S0(n5798), .S1(n5972), .Q(n436) );
  MUX41X1 U5487 ( .IN1(\FIFO[32][3] ), .IN3(\FIFO[34][3] ), .IN2(\FIFO[33][3] ), .IN4(\FIFO[35][3] ), .S0(n5798), .S1(n5895), .Q(n437) );
  MUX41X1 U5488 ( .IN1(n437), .IN3(n435), .IN2(n436), .IN4(n434), .S0(n5737), 
        .S1(n5780), .Q(n438) );
  MUX41X1 U5489 ( .IN1(\FIFO[28][3] ), .IN3(\FIFO[30][3] ), .IN2(\FIFO[29][3] ), .IN4(\FIFO[31][3] ), .S0(n5798), .S1(n5886), .Q(n439) );
  MUX41X1 U5490 ( .IN1(\FIFO[24][3] ), .IN3(\FIFO[26][3] ), .IN2(\FIFO[25][3] ), .IN4(\FIFO[27][3] ), .S0(n5798), .S1(n5875), .Q(n440) );
  MUX41X1 U5491 ( .IN1(\FIFO[20][3] ), .IN3(\FIFO[22][3] ), .IN2(\FIFO[21][3] ), .IN4(\FIFO[23][3] ), .S0(n5798), .S1(n5884), .Q(n441) );
  MUX41X1 U5492 ( .IN1(\FIFO[16][3] ), .IN3(\FIFO[18][3] ), .IN2(\FIFO[17][3] ), .IN4(\FIFO[19][3] ), .S0(n5798), .S1(n5885), .Q(n442) );
  MUX41X1 U5493 ( .IN1(n442), .IN3(n440), .IN2(n441), .IN4(n439), .S0(n5737), 
        .S1(N17), .Q(n443) );
  MUX41X1 U5494 ( .IN1(\FIFO[12][3] ), .IN3(\FIFO[14][3] ), .IN2(\FIFO[13][3] ), .IN4(\FIFO[15][3] ), .S0(n5799), .S1(n5895), .Q(n444) );
  MUX41X1 U5495 ( .IN1(\FIFO[8][3] ), .IN3(\FIFO[10][3] ), .IN2(\FIFO[9][3] ), 
        .IN4(\FIFO[11][3] ), .S0(n5799), .S1(n5882), .Q(n445) );
  MUX41X1 U5496 ( .IN1(\FIFO[4][3] ), .IN3(\FIFO[6][3] ), .IN2(\FIFO[5][3] ), 
        .IN4(\FIFO[7][3] ), .S0(n5799), .S1(n5967), .Q(n446) );
  MUX41X1 U5497 ( .IN1(\FIFO[0][3] ), .IN3(\FIFO[2][3] ), .IN2(\FIFO[1][3] ), 
        .IN4(\FIFO[3][3] ), .S0(n5799), .S1(n5968), .Q(n447) );
  MUX41X1 U5498 ( .IN1(n447), .IN3(n445), .IN2(n446), .IN4(n444), .S0(n5737), 
        .S1(n5780), .Q(n448) );
  MUX41X1 U5499 ( .IN1(n448), .IN3(n438), .IN2(n443), .IN4(n433), .S0(n5726), 
        .S1(n5730), .Q(n449) );
  MUX21X1 U5500 ( .IN1(n449), .IN2(n428), .S(N21), .Q(N247) );
  MUX41X1 U5501 ( .IN1(\FIFO[124][4] ), .IN3(\FIFO[126][4] ), .IN2(
        \FIFO[125][4] ), .IN4(\FIFO[127][4] ), .S0(n5799), .S1(n5893), .Q(n450) );
  MUX41X1 U5502 ( .IN1(\FIFO[120][4] ), .IN3(\FIFO[122][4] ), .IN2(
        \FIFO[121][4] ), .IN4(\FIFO[123][4] ), .S0(n5799), .S1(n5883), .Q(n451) );
  MUX41X1 U5503 ( .IN1(\FIFO[116][4] ), .IN3(\FIFO[118][4] ), .IN2(
        \FIFO[117][4] ), .IN4(\FIFO[119][4] ), .S0(n5799), .S1(n5880), .Q(n452) );
  MUX41X1 U5504 ( .IN1(\FIFO[112][4] ), .IN3(\FIFO[114][4] ), .IN2(
        \FIFO[113][4] ), .IN4(\FIFO[115][4] ), .S0(n5799), .S1(n5879), .Q(n453) );
  MUX41X1 U5505 ( .IN1(n453), .IN3(n451), .IN2(n452), .IN4(n450), .S0(n5737), 
        .S1(n5778), .Q(n454) );
  MUX41X1 U5506 ( .IN1(\FIFO[108][4] ), .IN3(\FIFO[110][4] ), .IN2(
        \FIFO[109][4] ), .IN4(\FIFO[111][4] ), .S0(n5799), .S1(n5881), .Q(n455) );
  MUX41X1 U5507 ( .IN1(\FIFO[104][4] ), .IN3(\FIFO[106][4] ), .IN2(
        \FIFO[105][4] ), .IN4(\FIFO[107][4] ), .S0(n5799), .S1(n5970), .Q(n456) );
  MUX41X1 U5508 ( .IN1(\FIFO[100][4] ), .IN3(\FIFO[102][4] ), .IN2(
        \FIFO[101][4] ), .IN4(\FIFO[103][4] ), .S0(n5799), .S1(n5894), .Q(n457) );
  MUX41X1 U5509 ( .IN1(\FIFO[96][4] ), .IN3(\FIFO[98][4] ), .IN2(\FIFO[97][4] ), .IN4(\FIFO[99][4] ), .S0(n5799), .S1(n5878), .Q(n458) );
  MUX41X1 U5510 ( .IN1(n458), .IN3(n456), .IN2(n457), .IN4(n455), .S0(n5737), 
        .S1(n5776), .Q(n459) );
  MUX41X1 U5511 ( .IN1(\FIFO[92][4] ), .IN3(\FIFO[94][4] ), .IN2(\FIFO[93][4] ), .IN4(\FIFO[95][4] ), .S0(n5800), .S1(n5886), .Q(n460) );
  MUX41X1 U5512 ( .IN1(\FIFO[88][4] ), .IN3(\FIFO[90][4] ), .IN2(\FIFO[89][4] ), .IN4(\FIFO[91][4] ), .S0(n5800), .S1(n5876), .Q(n461) );
  MUX41X1 U5513 ( .IN1(\FIFO[84][4] ), .IN3(\FIFO[86][4] ), .IN2(\FIFO[85][4] ), .IN4(\FIFO[87][4] ), .S0(n5800), .S1(n5965), .Q(n462) );
  MUX41X1 U5514 ( .IN1(\FIFO[80][4] ), .IN3(\FIFO[82][4] ), .IN2(\FIFO[81][4] ), .IN4(\FIFO[83][4] ), .S0(n5800), .S1(n5966), .Q(n463) );
  MUX41X1 U5515 ( .IN1(n463), .IN3(n461), .IN2(n462), .IN4(n460), .S0(n5737), 
        .S1(n5779), .Q(n465) );
  MUX41X1 U5516 ( .IN1(\FIFO[76][4] ), .IN3(\FIFO[78][4] ), .IN2(\FIFO[77][4] ), .IN4(\FIFO[79][4] ), .S0(n5800), .S1(n5875), .Q(n466) );
  MUX41X1 U5517 ( .IN1(\FIFO[72][4] ), .IN3(\FIFO[74][4] ), .IN2(\FIFO[73][4] ), .IN4(\FIFO[75][4] ), .S0(n5800), .S1(n5877), .Q(n4563) );
  MUX41X1 U5518 ( .IN1(\FIFO[68][4] ), .IN3(\FIFO[70][4] ), .IN2(\FIFO[69][4] ), .IN4(\FIFO[71][4] ), .S0(n5800), .S1(n5874), .Q(n4564) );
  MUX41X1 U5519 ( .IN1(\FIFO[64][4] ), .IN3(\FIFO[66][4] ), .IN2(\FIFO[65][4] ), .IN4(\FIFO[67][4] ), .S0(n5800), .S1(n5894), .Q(n4565) );
  MUX41X1 U5520 ( .IN1(n4565), .IN3(n4563), .IN2(n4564), .IN4(n466), .S0(n5737), .S1(n5777), .Q(n4566) );
  MUX41X1 U5521 ( .IN1(n4566), .IN3(n459), .IN2(n465), .IN4(n454), .S0(n5726), 
        .S1(n5730), .Q(n4567) );
  MUX41X1 U5522 ( .IN1(\FIFO[60][4] ), .IN3(\FIFO[62][4] ), .IN2(\FIFO[61][4] ), .IN4(\FIFO[63][4] ), .S0(n5800), .S1(n5893), .Q(n4568) );
  MUX41X1 U5523 ( .IN1(\FIFO[56][4] ), .IN3(\FIFO[58][4] ), .IN2(\FIFO[57][4] ), .IN4(\FIFO[59][4] ), .S0(n5800), .S1(n5896), .Q(n4569) );
  MUX41X1 U5524 ( .IN1(\FIFO[52][4] ), .IN3(\FIFO[54][4] ), .IN2(\FIFO[53][4] ), .IN4(\FIFO[55][4] ), .S0(n5800), .S1(n5969), .Q(n4570) );
  MUX41X1 U5525 ( .IN1(\FIFO[48][4] ), .IN3(\FIFO[50][4] ), .IN2(\FIFO[49][4] ), .IN4(\FIFO[51][4] ), .S0(n5800), .S1(n5970), .Q(n4571) );
  MUX41X1 U5526 ( .IN1(n4571), .IN3(n4569), .IN2(n4570), .IN4(n4568), .S0(
        n5737), .S1(n5777), .Q(n4572) );
  MUX41X1 U5527 ( .IN1(\FIFO[44][4] ), .IN3(\FIFO[46][4] ), .IN2(\FIFO[45][4] ), .IN4(\FIFO[47][4] ), .S0(n5801), .S1(n5891), .Q(n4573) );
  MUX41X1 U5528 ( .IN1(\FIFO[40][4] ), .IN3(\FIFO[42][4] ), .IN2(\FIFO[41][4] ), .IN4(\FIFO[43][4] ), .S0(n5801), .S1(n5892), .Q(n4574) );
  MUX41X1 U5529 ( .IN1(\FIFO[36][4] ), .IN3(\FIFO[38][4] ), .IN2(\FIFO[37][4] ), .IN4(\FIFO[39][4] ), .S0(n5801), .S1(n5971), .Q(n4575) );
  MUX41X1 U5530 ( .IN1(\FIFO[32][4] ), .IN3(\FIFO[34][4] ), .IN2(\FIFO[33][4] ), .IN4(\FIFO[35][4] ), .S0(n5801), .S1(n5972), .Q(n4576) );
  MUX41X1 U5531 ( .IN1(n4576), .IN3(n4574), .IN2(n4575), .IN4(n4573), .S0(
        n5737), .S1(n5781), .Q(n4577) );
  MUX41X1 U5532 ( .IN1(\FIFO[28][4] ), .IN3(\FIFO[30][4] ), .IN2(\FIFO[29][4] ), .IN4(\FIFO[31][4] ), .S0(n5801), .S1(n5888), .Q(n4578) );
  MUX41X1 U5533 ( .IN1(\FIFO[24][4] ), .IN3(\FIFO[26][4] ), .IN2(\FIFO[25][4] ), .IN4(\FIFO[27][4] ), .S0(n5801), .S1(n5874), .Q(n4579) );
  MUX41X1 U5534 ( .IN1(\FIFO[20][4] ), .IN3(\FIFO[22][4] ), .IN2(\FIFO[21][4] ), .IN4(\FIFO[23][4] ), .S0(n5801), .S1(n5886), .Q(n4580) );
  MUX41X1 U5535 ( .IN1(\FIFO[16][4] ), .IN3(\FIFO[18][4] ), .IN2(\FIFO[17][4] ), .IN4(\FIFO[19][4] ), .S0(n5801), .S1(n5887), .Q(n4581) );
  MUX41X1 U5536 ( .IN1(n4581), .IN3(n4579), .IN2(n4580), .IN4(n4578), .S0(
        n5737), .S1(N17), .Q(n4582) );
  MUX41X1 U5537 ( .IN1(\FIFO[12][4] ), .IN3(\FIFO[14][4] ), .IN2(\FIFO[13][4] ), .IN4(\FIFO[15][4] ), .S0(n5801), .S1(n5965), .Q(n4583) );
  MUX41X1 U5538 ( .IN1(\FIFO[8][4] ), .IN3(\FIFO[10][4] ), .IN2(\FIFO[9][4] ), 
        .IN4(\FIFO[11][4] ), .S0(n5801), .S1(n5890), .Q(n4584) );
  MUX41X1 U5539 ( .IN1(\FIFO[4][4] ), .IN3(\FIFO[6][4] ), .IN2(\FIFO[5][4] ), 
        .IN4(\FIFO[7][4] ), .S0(n5801), .S1(n5889), .Q(n4585) );
  MUX41X1 U5540 ( .IN1(\FIFO[0][4] ), .IN3(\FIFO[2][4] ), .IN2(\FIFO[1][4] ), 
        .IN4(\FIFO[3][4] ), .S0(n5801), .S1(n5972), .Q(n4586) );
  MUX41X1 U5541 ( .IN1(n4586), .IN3(n4584), .IN2(n4585), .IN4(n4583), .S0(
        n5737), .S1(n5781), .Q(n4587) );
  MUX41X1 U5542 ( .IN1(n4587), .IN3(n4577), .IN2(n4582), .IN4(n4572), .S0(
        n5726), .S1(n5730), .Q(n4588) );
  MUX21X1 U5543 ( .IN1(n4588), .IN2(n4567), .S(N21), .Q(N246) );
  MUX41X1 U5544 ( .IN1(\FIFO[124][5] ), .IN3(\FIFO[126][5] ), .IN2(
        \FIFO[125][5] ), .IN4(\FIFO[127][5] ), .S0(n5802), .S1(n5878), .Q(
        n4589) );
  MUX41X1 U5545 ( .IN1(\FIFO[120][5] ), .IN3(\FIFO[122][5] ), .IN2(
        \FIFO[121][5] ), .IN4(\FIFO[123][5] ), .S0(n5802), .S1(n5890), .Q(
        n4590) );
  MUX41X1 U5546 ( .IN1(\FIFO[116][5] ), .IN3(\FIFO[118][5] ), .IN2(
        \FIFO[117][5] ), .IN4(\FIFO[119][5] ), .S0(n5802), .S1(n5882), .Q(
        n4591) );
  MUX41X1 U5547 ( .IN1(\FIFO[112][5] ), .IN3(\FIFO[114][5] ), .IN2(
        \FIFO[113][5] ), .IN4(\FIFO[115][5] ), .S0(n5802), .S1(n5879), .Q(
        n4592) );
  MUX41X1 U5548 ( .IN1(n4592), .IN3(n4590), .IN2(n4591), .IN4(n4589), .S0(
        n5738), .S1(n5759), .Q(n4593) );
  MUX41X1 U5549 ( .IN1(\FIFO[108][5] ), .IN3(\FIFO[110][5] ), .IN2(
        \FIFO[109][5] ), .IN4(\FIFO[111][5] ), .S0(n5802), .S1(n5885), .Q(
        n4594) );
  MUX41X1 U5550 ( .IN1(\FIFO[104][5] ), .IN3(\FIFO[106][5] ), .IN2(
        \FIFO[105][5] ), .IN4(\FIFO[107][5] ), .S0(n5802), .S1(n5896), .Q(
        n4595) );
  MUX41X1 U5551 ( .IN1(\FIFO[100][5] ), .IN3(\FIFO[102][5] ), .IN2(
        \FIFO[101][5] ), .IN4(\FIFO[103][5] ), .S0(n5802), .S1(n5883), .Q(
        n4596) );
  MUX41X1 U5552 ( .IN1(\FIFO[96][5] ), .IN3(\FIFO[98][5] ), .IN2(\FIFO[97][5] ), .IN4(\FIFO[99][5] ), .S0(n5802), .S1(n5884), .Q(n4597) );
  MUX41X1 U5553 ( .IN1(n4597), .IN3(n4595), .IN2(n4596), .IN4(n4594), .S0(
        n5738), .S1(n5759), .Q(n4598) );
  MUX41X1 U5554 ( .IN1(\FIFO[92][5] ), .IN3(\FIFO[94][5] ), .IN2(\FIFO[93][5] ), .IN4(\FIFO[95][5] ), .S0(n5802), .S1(n5880), .Q(n4599) );
  MUX41X1 U5555 ( .IN1(\FIFO[88][5] ), .IN3(\FIFO[90][5] ), .IN2(\FIFO[89][5] ), .IN4(\FIFO[91][5] ), .S0(n5802), .S1(n5881), .Q(n4600) );
  MUX41X1 U5556 ( .IN1(\FIFO[84][5] ), .IN3(\FIFO[86][5] ), .IN2(\FIFO[85][5] ), .IN4(\FIFO[87][5] ), .S0(n5802), .S1(n5967), .Q(n4601) );
  MUX41X1 U5557 ( .IN1(\FIFO[80][5] ), .IN3(\FIFO[82][5] ), .IN2(\FIFO[81][5] ), .IN4(\FIFO[83][5] ), .S0(n5802), .S1(n5968), .Q(n4602) );
  MUX41X1 U5558 ( .IN1(n4602), .IN3(n4600), .IN2(n4601), .IN4(n4599), .S0(
        n5738), .S1(n5759), .Q(n4603) );
  MUX41X1 U5559 ( .IN1(\FIFO[76][5] ), .IN3(\FIFO[78][5] ), .IN2(\FIFO[77][5] ), .IN4(\FIFO[79][5] ), .S0(n5803), .S1(n5897), .Q(n4604) );
  MUX41X1 U5560 ( .IN1(\FIFO[72][5] ), .IN3(\FIFO[74][5] ), .IN2(\FIFO[73][5] ), .IN4(\FIFO[75][5] ), .S0(n5803), .S1(n5897), .Q(n4605) );
  MUX41X1 U5561 ( .IN1(\FIFO[68][5] ), .IN3(\FIFO[70][5] ), .IN2(\FIFO[69][5] ), .IN4(\FIFO[71][5] ), .S0(n5803), .S1(n5897), .Q(n4606) );
  MUX41X1 U5562 ( .IN1(\FIFO[64][5] ), .IN3(\FIFO[66][5] ), .IN2(\FIFO[65][5] ), .IN4(\FIFO[67][5] ), .S0(n5803), .S1(n5897), .Q(n4607) );
  MUX41X1 U5563 ( .IN1(n4607), .IN3(n4605), .IN2(n4606), .IN4(n4604), .S0(
        n5738), .S1(n5759), .Q(n4608) );
  MUX41X1 U5564 ( .IN1(n4608), .IN3(n4598), .IN2(n4603), .IN4(n4593), .S0(
        n5726), .S1(n5730), .Q(n4609) );
  MUX41X1 U5565 ( .IN1(\FIFO[60][5] ), .IN3(\FIFO[62][5] ), .IN2(\FIFO[61][5] ), .IN4(\FIFO[63][5] ), .S0(n5803), .S1(n5897), .Q(n4610) );
  MUX41X1 U5566 ( .IN1(\FIFO[56][5] ), .IN3(\FIFO[58][5] ), .IN2(\FIFO[57][5] ), .IN4(\FIFO[59][5] ), .S0(n5803), .S1(n5897), .Q(n4611) );
  MUX41X1 U5567 ( .IN1(\FIFO[52][5] ), .IN3(\FIFO[54][5] ), .IN2(\FIFO[53][5] ), .IN4(\FIFO[55][5] ), .S0(n5803), .S1(n5897), .Q(n4612) );
  MUX41X1 U5568 ( .IN1(\FIFO[48][5] ), .IN3(\FIFO[50][5] ), .IN2(\FIFO[49][5] ), .IN4(\FIFO[51][5] ), .S0(n5803), .S1(n5897), .Q(n4613) );
  MUX41X1 U5569 ( .IN1(n4613), .IN3(n4611), .IN2(n4612), .IN4(n4610), .S0(
        n5738), .S1(n5759), .Q(n4614) );
  MUX41X1 U5570 ( .IN1(\FIFO[44][5] ), .IN3(\FIFO[46][5] ), .IN2(\FIFO[45][5] ), .IN4(\FIFO[47][5] ), .S0(n5803), .S1(n5897), .Q(n4615) );
  MUX41X1 U5571 ( .IN1(\FIFO[40][5] ), .IN3(\FIFO[42][5] ), .IN2(\FIFO[41][5] ), .IN4(\FIFO[43][5] ), .S0(n5803), .S1(n5897), .Q(n4616) );
  MUX41X1 U5572 ( .IN1(\FIFO[36][5] ), .IN3(\FIFO[38][5] ), .IN2(\FIFO[37][5] ), .IN4(\FIFO[39][5] ), .S0(n5803), .S1(n5897), .Q(n4617) );
  MUX41X1 U5573 ( .IN1(\FIFO[32][5] ), .IN3(\FIFO[34][5] ), .IN2(\FIFO[33][5] ), .IN4(\FIFO[35][5] ), .S0(n5803), .S1(n5897), .Q(n4618) );
  MUX41X1 U5574 ( .IN1(n4618), .IN3(n4616), .IN2(n4617), .IN4(n4615), .S0(
        n5738), .S1(n5759), .Q(n4619) );
  MUX41X1 U5575 ( .IN1(\FIFO[28][5] ), .IN3(\FIFO[30][5] ), .IN2(\FIFO[29][5] ), .IN4(\FIFO[31][5] ), .S0(n5804), .S1(n5898), .Q(n4620) );
  MUX41X1 U5576 ( .IN1(\FIFO[24][5] ), .IN3(\FIFO[26][5] ), .IN2(\FIFO[25][5] ), .IN4(\FIFO[27][5] ), .S0(n5804), .S1(n5898), .Q(n4621) );
  MUX41X1 U5577 ( .IN1(\FIFO[20][5] ), .IN3(\FIFO[22][5] ), .IN2(\FIFO[21][5] ), .IN4(\FIFO[23][5] ), .S0(n5804), .S1(n5898), .Q(n4622) );
  MUX41X1 U5578 ( .IN1(\FIFO[16][5] ), .IN3(\FIFO[18][5] ), .IN2(\FIFO[17][5] ), .IN4(\FIFO[19][5] ), .S0(n5804), .S1(n5898), .Q(n4623) );
  MUX41X1 U5579 ( .IN1(n4623), .IN3(n4621), .IN2(n4622), .IN4(n4620), .S0(
        n5738), .S1(n5759), .Q(n4624) );
  MUX41X1 U5580 ( .IN1(\FIFO[12][5] ), .IN3(\FIFO[14][5] ), .IN2(\FIFO[13][5] ), .IN4(\FIFO[15][5] ), .S0(n5804), .S1(n5898), .Q(n4625) );
  MUX41X1 U5581 ( .IN1(\FIFO[8][5] ), .IN3(\FIFO[10][5] ), .IN2(\FIFO[9][5] ), 
        .IN4(\FIFO[11][5] ), .S0(n5804), .S1(n5898), .Q(n4626) );
  MUX41X1 U5582 ( .IN1(\FIFO[4][5] ), .IN3(\FIFO[6][5] ), .IN2(\FIFO[5][5] ), 
        .IN4(\FIFO[7][5] ), .S0(n5804), .S1(n5898), .Q(n4627) );
  MUX41X1 U5583 ( .IN1(\FIFO[0][5] ), .IN3(\FIFO[2][5] ), .IN2(\FIFO[1][5] ), 
        .IN4(\FIFO[3][5] ), .S0(n5804), .S1(n5898), .Q(n4628) );
  MUX41X1 U5584 ( .IN1(n4628), .IN3(n4626), .IN2(n4627), .IN4(n4625), .S0(
        n5738), .S1(n5759), .Q(n4629) );
  MUX41X1 U5585 ( .IN1(n4629), .IN3(n4619), .IN2(n4624), .IN4(n4614), .S0(
        n5726), .S1(n5730), .Q(n4630) );
  MUX21X1 U5586 ( .IN1(n4630), .IN2(n4609), .S(N21), .Q(N245) );
  MUX41X1 U5587 ( .IN1(\FIFO[124][6] ), .IN3(\FIFO[126][6] ), .IN2(
        \FIFO[125][6] ), .IN4(\FIFO[127][6] ), .S0(n5804), .S1(n5898), .Q(
        n4631) );
  MUX41X1 U5588 ( .IN1(\FIFO[120][6] ), .IN3(\FIFO[122][6] ), .IN2(
        \FIFO[121][6] ), .IN4(\FIFO[123][6] ), .S0(n5804), .S1(n5898), .Q(
        n4632) );
  MUX41X1 U5589 ( .IN1(\FIFO[116][6] ), .IN3(\FIFO[118][6] ), .IN2(
        \FIFO[117][6] ), .IN4(\FIFO[119][6] ), .S0(n5804), .S1(n5898), .Q(
        n4633) );
  MUX41X1 U5590 ( .IN1(\FIFO[112][6] ), .IN3(\FIFO[114][6] ), .IN2(
        \FIFO[113][6] ), .IN4(\FIFO[115][6] ), .S0(n5804), .S1(n5898), .Q(
        n4634) );
  MUX41X1 U5591 ( .IN1(n4634), .IN3(n4632), .IN2(n4633), .IN4(n4631), .S0(
        n5738), .S1(n5759), .Q(n4635) );
  MUX41X1 U5592 ( .IN1(\FIFO[108][6] ), .IN3(\FIFO[110][6] ), .IN2(
        \FIFO[109][6] ), .IN4(\FIFO[111][6] ), .S0(n5805), .S1(n5899), .Q(
        n4636) );
  MUX41X1 U5593 ( .IN1(\FIFO[104][6] ), .IN3(\FIFO[106][6] ), .IN2(
        \FIFO[105][6] ), .IN4(\FIFO[107][6] ), .S0(n5805), .S1(n5899), .Q(
        n4637) );
  MUX41X1 U5594 ( .IN1(\FIFO[100][6] ), .IN3(\FIFO[102][6] ), .IN2(
        \FIFO[101][6] ), .IN4(\FIFO[103][6] ), .S0(n5805), .S1(n5899), .Q(
        n4638) );
  MUX41X1 U5595 ( .IN1(\FIFO[96][6] ), .IN3(\FIFO[98][6] ), .IN2(\FIFO[97][6] ), .IN4(\FIFO[99][6] ), .S0(n5805), .S1(n5899), .Q(n4639) );
  MUX41X1 U5596 ( .IN1(n4639), .IN3(n4637), .IN2(n4638), .IN4(n4636), .S0(
        n5738), .S1(n5759), .Q(n4640) );
  MUX41X1 U5597 ( .IN1(\FIFO[92][6] ), .IN3(\FIFO[94][6] ), .IN2(\FIFO[93][6] ), .IN4(\FIFO[95][6] ), .S0(n5805), .S1(n5899), .Q(n4641) );
  MUX41X1 U5598 ( .IN1(\FIFO[88][6] ), .IN3(\FIFO[90][6] ), .IN2(\FIFO[89][6] ), .IN4(\FIFO[91][6] ), .S0(n5805), .S1(n5899), .Q(n4642) );
  MUX41X1 U5599 ( .IN1(\FIFO[84][6] ), .IN3(\FIFO[86][6] ), .IN2(\FIFO[85][6] ), .IN4(\FIFO[87][6] ), .S0(n5805), .S1(n5899), .Q(n4643) );
  MUX41X1 U5600 ( .IN1(\FIFO[80][6] ), .IN3(\FIFO[82][6] ), .IN2(\FIFO[81][6] ), .IN4(\FIFO[83][6] ), .S0(n5805), .S1(n5899), .Q(n4644) );
  MUX41X1 U5601 ( .IN1(n4644), .IN3(n4642), .IN2(n4643), .IN4(n4641), .S0(
        n5738), .S1(n5759), .Q(n4645) );
  MUX41X1 U5602 ( .IN1(\FIFO[76][6] ), .IN3(\FIFO[78][6] ), .IN2(\FIFO[77][6] ), .IN4(\FIFO[79][6] ), .S0(n5805), .S1(n5899), .Q(n4646) );
  MUX41X1 U5603 ( .IN1(\FIFO[72][6] ), .IN3(\FIFO[74][6] ), .IN2(\FIFO[73][6] ), .IN4(\FIFO[75][6] ), .S0(n5805), .S1(n5899), .Q(n4647) );
  MUX41X1 U5604 ( .IN1(\FIFO[68][6] ), .IN3(\FIFO[70][6] ), .IN2(\FIFO[69][6] ), .IN4(\FIFO[71][6] ), .S0(n5805), .S1(n5899), .Q(n4648) );
  MUX41X1 U5605 ( .IN1(\FIFO[64][6] ), .IN3(\FIFO[66][6] ), .IN2(\FIFO[65][6] ), .IN4(\FIFO[67][6] ), .S0(n5805), .S1(n5899), .Q(n4649) );
  MUX41X1 U5606 ( .IN1(n4649), .IN3(n4647), .IN2(n4648), .IN4(n4646), .S0(
        n5738), .S1(n5759), .Q(n4650) );
  MUX41X1 U5607 ( .IN1(n4650), .IN3(n4640), .IN2(n4645), .IN4(n4635), .S0(
        n5726), .S1(n5730), .Q(n4651) );
  MUX41X1 U5608 ( .IN1(\FIFO[60][6] ), .IN3(\FIFO[62][6] ), .IN2(\FIFO[61][6] ), .IN4(\FIFO[63][6] ), .S0(n5806), .S1(n5900), .Q(n4652) );
  MUX41X1 U5609 ( .IN1(\FIFO[56][6] ), .IN3(\FIFO[58][6] ), .IN2(\FIFO[57][6] ), .IN4(\FIFO[59][6] ), .S0(n5806), .S1(n5900), .Q(n4653) );
  MUX41X1 U5610 ( .IN1(\FIFO[52][6] ), .IN3(\FIFO[54][6] ), .IN2(\FIFO[53][6] ), .IN4(\FIFO[55][6] ), .S0(n5806), .S1(n5900), .Q(n4654) );
  MUX41X1 U5611 ( .IN1(\FIFO[48][6] ), .IN3(\FIFO[50][6] ), .IN2(\FIFO[49][6] ), .IN4(\FIFO[51][6] ), .S0(n5806), .S1(n5900), .Q(n4655) );
  MUX41X1 U5612 ( .IN1(n4655), .IN3(n4653), .IN2(n4654), .IN4(n4652), .S0(
        n5739), .S1(n5775), .Q(n4656) );
  MUX41X1 U5613 ( .IN1(\FIFO[44][6] ), .IN3(\FIFO[46][6] ), .IN2(\FIFO[45][6] ), .IN4(\FIFO[47][6] ), .S0(n5806), .S1(n5900), .Q(n4657) );
  MUX41X1 U5614 ( .IN1(\FIFO[40][6] ), .IN3(\FIFO[42][6] ), .IN2(\FIFO[41][6] ), .IN4(\FIFO[43][6] ), .S0(n5806), .S1(n5900), .Q(n4658) );
  MUX41X1 U5615 ( .IN1(\FIFO[36][6] ), .IN3(\FIFO[38][6] ), .IN2(\FIFO[37][6] ), .IN4(\FIFO[39][6] ), .S0(n5806), .S1(n5900), .Q(n4659) );
  MUX41X1 U5616 ( .IN1(\FIFO[32][6] ), .IN3(\FIFO[34][6] ), .IN2(\FIFO[33][6] ), .IN4(\FIFO[35][6] ), .S0(n5806), .S1(n5900), .Q(n4660) );
  MUX41X1 U5617 ( .IN1(n4660), .IN3(n4658), .IN2(n4659), .IN4(n4657), .S0(
        n5739), .S1(n5775), .Q(n4661) );
  MUX41X1 U5618 ( .IN1(\FIFO[28][6] ), .IN3(\FIFO[30][6] ), .IN2(\FIFO[29][6] ), .IN4(\FIFO[31][6] ), .S0(n5806), .S1(n5900), .Q(n4662) );
  MUX41X1 U5619 ( .IN1(\FIFO[24][6] ), .IN3(\FIFO[26][6] ), .IN2(\FIFO[25][6] ), .IN4(\FIFO[27][6] ), .S0(n5806), .S1(n5900), .Q(n4663) );
  MUX41X1 U5620 ( .IN1(\FIFO[20][6] ), .IN3(\FIFO[22][6] ), .IN2(\FIFO[21][6] ), .IN4(\FIFO[23][6] ), .S0(n5806), .S1(n5900), .Q(n4664) );
  MUX41X1 U5621 ( .IN1(\FIFO[16][6] ), .IN3(\FIFO[18][6] ), .IN2(\FIFO[17][6] ), .IN4(\FIFO[19][6] ), .S0(n5806), .S1(n5900), .Q(n4665) );
  MUX41X1 U5622 ( .IN1(n4665), .IN3(n4663), .IN2(n4664), .IN4(n4662), .S0(
        n5739), .S1(n5758), .Q(n4666) );
  MUX41X1 U5623 ( .IN1(\FIFO[12][6] ), .IN3(\FIFO[14][6] ), .IN2(\FIFO[13][6] ), .IN4(\FIFO[15][6] ), .S0(n5807), .S1(n5901), .Q(n4667) );
  MUX41X1 U5624 ( .IN1(\FIFO[8][6] ), .IN3(\FIFO[10][6] ), .IN2(\FIFO[9][6] ), 
        .IN4(\FIFO[11][6] ), .S0(n5807), .S1(n5901), .Q(n4668) );
  MUX41X1 U5625 ( .IN1(\FIFO[4][6] ), .IN3(\FIFO[6][6] ), .IN2(\FIFO[5][6] ), 
        .IN4(\FIFO[7][6] ), .S0(n5807), .S1(n5901), .Q(n4669) );
  MUX41X1 U5626 ( .IN1(\FIFO[0][6] ), .IN3(\FIFO[2][6] ), .IN2(\FIFO[1][6] ), 
        .IN4(\FIFO[3][6] ), .S0(n5807), .S1(n5901), .Q(n4670) );
  MUX41X1 U5627 ( .IN1(n4670), .IN3(n4668), .IN2(n4669), .IN4(n4667), .S0(
        n5739), .S1(n5758), .Q(n4671) );
  MUX41X1 U5628 ( .IN1(n4671), .IN3(n4661), .IN2(n4666), .IN4(n4656), .S0(
        n5726), .S1(n5730), .Q(n4672) );
  MUX21X1 U5629 ( .IN1(n4672), .IN2(n4651), .S(N21), .Q(N244) );
  MUX41X1 U5630 ( .IN1(\FIFO[124][7] ), .IN3(\FIFO[126][7] ), .IN2(
        \FIFO[125][7] ), .IN4(\FIFO[127][7] ), .S0(n5807), .S1(n5901), .Q(
        n4673) );
  MUX41X1 U5631 ( .IN1(\FIFO[120][7] ), .IN3(\FIFO[122][7] ), .IN2(
        \FIFO[121][7] ), .IN4(\FIFO[123][7] ), .S0(n5807), .S1(n5901), .Q(
        n4674) );
  MUX41X1 U5632 ( .IN1(\FIFO[116][7] ), .IN3(\FIFO[118][7] ), .IN2(
        \FIFO[117][7] ), .IN4(\FIFO[119][7] ), .S0(n5807), .S1(n5901), .Q(
        n4675) );
  MUX41X1 U5633 ( .IN1(\FIFO[112][7] ), .IN3(\FIFO[114][7] ), .IN2(
        \FIFO[113][7] ), .IN4(\FIFO[115][7] ), .S0(n5807), .S1(n5901), .Q(
        n4676) );
  MUX41X1 U5634 ( .IN1(n4676), .IN3(n4674), .IN2(n4675), .IN4(n4673), .S0(
        n5739), .S1(n5775), .Q(n4677) );
  MUX41X1 U5635 ( .IN1(\FIFO[108][7] ), .IN3(\FIFO[110][7] ), .IN2(
        \FIFO[109][7] ), .IN4(\FIFO[111][7] ), .S0(n5807), .S1(n5901), .Q(
        n4678) );
  MUX41X1 U5636 ( .IN1(\FIFO[104][7] ), .IN3(\FIFO[106][7] ), .IN2(
        \FIFO[105][7] ), .IN4(\FIFO[107][7] ), .S0(n5807), .S1(n5901), .Q(
        n4679) );
  MUX41X1 U5637 ( .IN1(\FIFO[100][7] ), .IN3(\FIFO[102][7] ), .IN2(
        \FIFO[101][7] ), .IN4(\FIFO[103][7] ), .S0(n5807), .S1(n5901), .Q(
        n4680) );
  MUX41X1 U5638 ( .IN1(\FIFO[96][7] ), .IN3(\FIFO[98][7] ), .IN2(\FIFO[97][7] ), .IN4(\FIFO[99][7] ), .S0(n5807), .S1(n5901), .Q(n4681) );
  MUX41X1 U5639 ( .IN1(n4681), .IN3(n4679), .IN2(n4680), .IN4(n4678), .S0(
        n5739), .S1(n5775), .Q(n4682) );
  MUX41X1 U5640 ( .IN1(\FIFO[92][7] ), .IN3(\FIFO[94][7] ), .IN2(\FIFO[93][7] ), .IN4(\FIFO[95][7] ), .S0(n5808), .S1(n5902), .Q(n4683) );
  MUX41X1 U5641 ( .IN1(\FIFO[88][7] ), .IN3(\FIFO[90][7] ), .IN2(\FIFO[89][7] ), .IN4(\FIFO[91][7] ), .S0(n5808), .S1(n5902), .Q(n4684) );
  MUX41X1 U5642 ( .IN1(\FIFO[84][7] ), .IN3(\FIFO[86][7] ), .IN2(\FIFO[85][7] ), .IN4(\FIFO[87][7] ), .S0(n5808), .S1(n5902), .Q(n4685) );
  MUX41X1 U5643 ( .IN1(\FIFO[80][7] ), .IN3(\FIFO[82][7] ), .IN2(\FIFO[81][7] ), .IN4(\FIFO[83][7] ), .S0(n5808), .S1(n5902), .Q(n4686) );
  MUX41X1 U5644 ( .IN1(n4686), .IN3(n4684), .IN2(n4685), .IN4(n4683), .S0(
        n5739), .S1(n5775), .Q(n4687) );
  MUX41X1 U5645 ( .IN1(\FIFO[76][7] ), .IN3(\FIFO[78][7] ), .IN2(\FIFO[77][7] ), .IN4(\FIFO[79][7] ), .S0(n5808), .S1(n5902), .Q(n4688) );
  MUX41X1 U5646 ( .IN1(\FIFO[72][7] ), .IN3(\FIFO[74][7] ), .IN2(\FIFO[73][7] ), .IN4(\FIFO[75][7] ), .S0(n5808), .S1(n5902), .Q(n4689) );
  MUX41X1 U5647 ( .IN1(\FIFO[68][7] ), .IN3(\FIFO[70][7] ), .IN2(\FIFO[69][7] ), .IN4(\FIFO[71][7] ), .S0(n5808), .S1(n5902), .Q(n4690) );
  MUX41X1 U5648 ( .IN1(\FIFO[64][7] ), .IN3(\FIFO[66][7] ), .IN2(\FIFO[65][7] ), .IN4(\FIFO[67][7] ), .S0(n5808), .S1(n5902), .Q(n4691) );
  MUX41X1 U5649 ( .IN1(n4691), .IN3(n4689), .IN2(n4690), .IN4(n4688), .S0(
        n5739), .S1(n5775), .Q(n4692) );
  MUX41X1 U5650 ( .IN1(n4692), .IN3(n4682), .IN2(n4687), .IN4(n4677), .S0(
        n5726), .S1(n5730), .Q(n4693) );
  MUX41X1 U5651 ( .IN1(\FIFO[60][7] ), .IN3(\FIFO[62][7] ), .IN2(\FIFO[61][7] ), .IN4(\FIFO[63][7] ), .S0(n5808), .S1(n5902), .Q(n4694) );
  MUX41X1 U5652 ( .IN1(\FIFO[56][7] ), .IN3(\FIFO[58][7] ), .IN2(\FIFO[57][7] ), .IN4(\FIFO[59][7] ), .S0(n5808), .S1(n5902), .Q(n4695) );
  MUX41X1 U5653 ( .IN1(\FIFO[52][7] ), .IN3(\FIFO[54][7] ), .IN2(\FIFO[53][7] ), .IN4(\FIFO[55][7] ), .S0(n5808), .S1(n5902), .Q(n4696) );
  MUX41X1 U5654 ( .IN1(\FIFO[48][7] ), .IN3(\FIFO[50][7] ), .IN2(\FIFO[49][7] ), .IN4(\FIFO[51][7] ), .S0(n5808), .S1(n5902), .Q(n4697) );
  MUX41X1 U5655 ( .IN1(n4697), .IN3(n4695), .IN2(n4696), .IN4(n4694), .S0(
        n5739), .S1(n5775), .Q(n4698) );
  MUX41X1 U5656 ( .IN1(\FIFO[44][7] ), .IN3(\FIFO[46][7] ), .IN2(\FIFO[45][7] ), .IN4(\FIFO[47][7] ), .S0(n5809), .S1(n5903), .Q(n4699) );
  MUX41X1 U5657 ( .IN1(\FIFO[40][7] ), .IN3(\FIFO[42][7] ), .IN2(\FIFO[41][7] ), .IN4(\FIFO[43][7] ), .S0(n5809), .S1(n5903), .Q(n4700) );
  MUX41X1 U5658 ( .IN1(\FIFO[36][7] ), .IN3(\FIFO[38][7] ), .IN2(\FIFO[37][7] ), .IN4(\FIFO[39][7] ), .S0(n5809), .S1(n5903), .Q(n4701) );
  MUX41X1 U5659 ( .IN1(\FIFO[32][7] ), .IN3(\FIFO[34][7] ), .IN2(\FIFO[33][7] ), .IN4(\FIFO[35][7] ), .S0(n5809), .S1(n5903), .Q(n4702) );
  MUX41X1 U5660 ( .IN1(n4702), .IN3(n4700), .IN2(n4701), .IN4(n4699), .S0(
        n5739), .S1(n5775), .Q(n4703) );
  MUX41X1 U5661 ( .IN1(\FIFO[28][7] ), .IN3(\FIFO[30][7] ), .IN2(\FIFO[29][7] ), .IN4(\FIFO[31][7] ), .S0(n5809), .S1(n5903), .Q(n4704) );
  MUX41X1 U5662 ( .IN1(\FIFO[24][7] ), .IN3(\FIFO[26][7] ), .IN2(\FIFO[25][7] ), .IN4(\FIFO[27][7] ), .S0(n5809), .S1(n5903), .Q(n4705) );
  MUX41X1 U5663 ( .IN1(\FIFO[20][7] ), .IN3(\FIFO[22][7] ), .IN2(\FIFO[21][7] ), .IN4(\FIFO[23][7] ), .S0(n5809), .S1(n5903), .Q(n4706) );
  MUX41X1 U5664 ( .IN1(\FIFO[16][7] ), .IN3(\FIFO[18][7] ), .IN2(\FIFO[17][7] ), .IN4(\FIFO[19][7] ), .S0(n5809), .S1(n5903), .Q(n4707) );
  MUX41X1 U5665 ( .IN1(n4707), .IN3(n4705), .IN2(n4706), .IN4(n4704), .S0(
        n5739), .S1(n5758), .Q(n4708) );
  MUX41X1 U5666 ( .IN1(\FIFO[12][7] ), .IN3(\FIFO[14][7] ), .IN2(\FIFO[13][7] ), .IN4(\FIFO[15][7] ), .S0(n5809), .S1(n5903), .Q(n4709) );
  MUX41X1 U5667 ( .IN1(\FIFO[8][7] ), .IN3(\FIFO[10][7] ), .IN2(\FIFO[9][7] ), 
        .IN4(\FIFO[11][7] ), .S0(n5809), .S1(n5903), .Q(n4710) );
  MUX41X1 U5668 ( .IN1(\FIFO[4][7] ), .IN3(\FIFO[6][7] ), .IN2(\FIFO[5][7] ), 
        .IN4(\FIFO[7][7] ), .S0(n5809), .S1(n5903), .Q(n4711) );
  MUX41X1 U5669 ( .IN1(\FIFO[0][7] ), .IN3(\FIFO[2][7] ), .IN2(\FIFO[1][7] ), 
        .IN4(\FIFO[3][7] ), .S0(n5809), .S1(n5903), .Q(n4712) );
  MUX41X1 U5670 ( .IN1(n4712), .IN3(n4710), .IN2(n4711), .IN4(n4709), .S0(
        n5739), .S1(n5758), .Q(n4713) );
  MUX41X1 U5671 ( .IN1(n4713), .IN3(n4703), .IN2(n4708), .IN4(n4698), .S0(
        n5726), .S1(n5730), .Q(n4714) );
  MUX21X1 U5672 ( .IN1(n4714), .IN2(n4693), .S(N21), .Q(N243) );
  MUX41X1 U5673 ( .IN1(\FIFO[124][8] ), .IN3(\FIFO[126][8] ), .IN2(
        \FIFO[125][8] ), .IN4(\FIFO[127][8] ), .S0(n5810), .S1(n5904), .Q(
        n4715) );
  MUX41X1 U5674 ( .IN1(\FIFO[120][8] ), .IN3(\FIFO[122][8] ), .IN2(
        \FIFO[121][8] ), .IN4(\FIFO[123][8] ), .S0(n5810), .S1(n5904), .Q(
        n4716) );
  MUX41X1 U5675 ( .IN1(\FIFO[116][8] ), .IN3(\FIFO[118][8] ), .IN2(
        \FIFO[117][8] ), .IN4(\FIFO[119][8] ), .S0(n5810), .S1(n5904), .Q(
        n4717) );
  MUX41X1 U5676 ( .IN1(\FIFO[112][8] ), .IN3(\FIFO[114][8] ), .IN2(
        \FIFO[113][8] ), .IN4(\FIFO[115][8] ), .S0(n5810), .S1(n5904), .Q(
        n4718) );
  MUX41X1 U5677 ( .IN1(n4718), .IN3(n4716), .IN2(n4717), .IN4(n4715), .S0(
        n5740), .S1(n5776), .Q(n4719) );
  MUX41X1 U5678 ( .IN1(\FIFO[108][8] ), .IN3(\FIFO[110][8] ), .IN2(
        \FIFO[109][8] ), .IN4(\FIFO[111][8] ), .S0(n5810), .S1(n5904), .Q(
        n4720) );
  MUX41X1 U5679 ( .IN1(\FIFO[104][8] ), .IN3(\FIFO[106][8] ), .IN2(
        \FIFO[105][8] ), .IN4(\FIFO[107][8] ), .S0(n5810), .S1(n5904), .Q(
        n4721) );
  MUX41X1 U5680 ( .IN1(\FIFO[100][8] ), .IN3(\FIFO[102][8] ), .IN2(
        \FIFO[101][8] ), .IN4(\FIFO[103][8] ), .S0(n5810), .S1(n5904), .Q(
        n4722) );
  MUX41X1 U5681 ( .IN1(\FIFO[96][8] ), .IN3(\FIFO[98][8] ), .IN2(\FIFO[97][8] ), .IN4(\FIFO[99][8] ), .S0(n5810), .S1(n5904), .Q(n4723) );
  MUX41X1 U5682 ( .IN1(n4723), .IN3(n4721), .IN2(n4722), .IN4(n4720), .S0(
        n5740), .S1(n5780), .Q(n4724) );
  MUX41X1 U5683 ( .IN1(\FIFO[92][8] ), .IN3(\FIFO[94][8] ), .IN2(\FIFO[93][8] ), .IN4(\FIFO[95][8] ), .S0(n5810), .S1(n5904), .Q(n4725) );
  MUX41X1 U5684 ( .IN1(\FIFO[88][8] ), .IN3(\FIFO[90][8] ), .IN2(\FIFO[89][8] ), .IN4(\FIFO[91][8] ), .S0(n5810), .S1(n5904), .Q(n4726) );
  MUX41X1 U5685 ( .IN1(\FIFO[84][8] ), .IN3(\FIFO[86][8] ), .IN2(\FIFO[85][8] ), .IN4(\FIFO[87][8] ), .S0(n5810), .S1(n5904), .Q(n4727) );
  MUX41X1 U5686 ( .IN1(\FIFO[80][8] ), .IN3(\FIFO[82][8] ), .IN2(\FIFO[81][8] ), .IN4(\FIFO[83][8] ), .S0(n5810), .S1(n5904), .Q(n4728) );
  MUX41X1 U5687 ( .IN1(n4728), .IN3(n4726), .IN2(n4727), .IN4(n4725), .S0(
        n5740), .S1(n5781), .Q(n4729) );
  MUX41X1 U5688 ( .IN1(\FIFO[76][8] ), .IN3(\FIFO[78][8] ), .IN2(\FIFO[77][8] ), .IN4(\FIFO[79][8] ), .S0(n5811), .S1(n5905), .Q(n4730) );
  MUX41X1 U5689 ( .IN1(\FIFO[72][8] ), .IN3(\FIFO[74][8] ), .IN2(\FIFO[73][8] ), .IN4(\FIFO[75][8] ), .S0(n5811), .S1(n5905), .Q(n4731) );
  MUX41X1 U5690 ( .IN1(\FIFO[68][8] ), .IN3(\FIFO[70][8] ), .IN2(\FIFO[69][8] ), .IN4(\FIFO[71][8] ), .S0(n5811), .S1(n5905), .Q(n4732) );
  MUX41X1 U5691 ( .IN1(\FIFO[64][8] ), .IN3(\FIFO[66][8] ), .IN2(\FIFO[65][8] ), .IN4(\FIFO[67][8] ), .S0(n5811), .S1(n5905), .Q(n4733) );
  MUX41X1 U5692 ( .IN1(n4733), .IN3(n4731), .IN2(n4732), .IN4(n4730), .S0(
        n5740), .S1(n5777), .Q(n4734) );
  MUX41X1 U5693 ( .IN1(n4734), .IN3(n4724), .IN2(n4729), .IN4(n4719), .S0(
        n5727), .S1(n5731), .Q(n4735) );
  MUX41X1 U5694 ( .IN1(\FIFO[60][8] ), .IN3(\FIFO[62][8] ), .IN2(\FIFO[61][8] ), .IN4(\FIFO[63][8] ), .S0(n5811), .S1(n5905), .Q(n4736) );
  MUX41X1 U5695 ( .IN1(\FIFO[56][8] ), .IN3(\FIFO[58][8] ), .IN2(\FIFO[57][8] ), .IN4(\FIFO[59][8] ), .S0(n5811), .S1(n5905), .Q(n4737) );
  MUX41X1 U5696 ( .IN1(\FIFO[52][8] ), .IN3(\FIFO[54][8] ), .IN2(\FIFO[53][8] ), .IN4(\FIFO[55][8] ), .S0(n5811), .S1(n5905), .Q(n4738) );
  MUX41X1 U5697 ( .IN1(\FIFO[48][8] ), .IN3(\FIFO[50][8] ), .IN2(\FIFO[49][8] ), .IN4(\FIFO[51][8] ), .S0(n5811), .S1(n5905), .Q(n4739) );
  MUX41X1 U5698 ( .IN1(n4739), .IN3(n4737), .IN2(n4738), .IN4(n4736), .S0(
        n5740), .S1(n5776), .Q(n4740) );
  MUX41X1 U5699 ( .IN1(\FIFO[44][8] ), .IN3(\FIFO[46][8] ), .IN2(\FIFO[45][8] ), .IN4(\FIFO[47][8] ), .S0(n5811), .S1(n5905), .Q(n4741) );
  MUX41X1 U5700 ( .IN1(\FIFO[40][8] ), .IN3(\FIFO[42][8] ), .IN2(\FIFO[41][8] ), .IN4(\FIFO[43][8] ), .S0(n5811), .S1(n5905), .Q(n4742) );
  MUX41X1 U5701 ( .IN1(\FIFO[36][8] ), .IN3(\FIFO[38][8] ), .IN2(\FIFO[37][8] ), .IN4(\FIFO[39][8] ), .S0(n5811), .S1(n5905), .Q(n4743) );
  MUX41X1 U5702 ( .IN1(\FIFO[32][8] ), .IN3(\FIFO[34][8] ), .IN2(\FIFO[33][8] ), .IN4(\FIFO[35][8] ), .S0(n5811), .S1(n5905), .Q(n4744) );
  MUX41X1 U5703 ( .IN1(n4744), .IN3(n4742), .IN2(n4743), .IN4(n4741), .S0(
        n5740), .S1(n5780), .Q(n4745) );
  MUX41X1 U5704 ( .IN1(\FIFO[28][8] ), .IN3(\FIFO[30][8] ), .IN2(\FIFO[29][8] ), .IN4(\FIFO[31][8] ), .S0(n5812), .S1(n5906), .Q(n4746) );
  MUX41X1 U5705 ( .IN1(\FIFO[24][8] ), .IN3(\FIFO[26][8] ), .IN2(\FIFO[25][8] ), .IN4(\FIFO[27][8] ), .S0(n5812), .S1(n5906), .Q(n4747) );
  MUX41X1 U5706 ( .IN1(\FIFO[20][8] ), .IN3(\FIFO[22][8] ), .IN2(\FIFO[21][8] ), .IN4(\FIFO[23][8] ), .S0(n5812), .S1(n5906), .Q(n4748) );
  MUX41X1 U5707 ( .IN1(\FIFO[16][8] ), .IN3(\FIFO[18][8] ), .IN2(\FIFO[17][8] ), .IN4(\FIFO[19][8] ), .S0(n5812), .S1(n5906), .Q(n4749) );
  MUX41X1 U5708 ( .IN1(n4749), .IN3(n4747), .IN2(n4748), .IN4(n4746), .S0(
        n5740), .S1(n5777), .Q(n4750) );
  MUX41X1 U5709 ( .IN1(\FIFO[12][8] ), .IN3(\FIFO[14][8] ), .IN2(\FIFO[13][8] ), .IN4(\FIFO[15][8] ), .S0(n5812), .S1(n5906), .Q(n4751) );
  MUX41X1 U5710 ( .IN1(\FIFO[8][8] ), .IN3(\FIFO[10][8] ), .IN2(\FIFO[9][8] ), 
        .IN4(\FIFO[11][8] ), .S0(n5812), .S1(n5906), .Q(n4752) );
  MUX41X1 U5711 ( .IN1(\FIFO[4][8] ), .IN3(\FIFO[6][8] ), .IN2(\FIFO[5][8] ), 
        .IN4(\FIFO[7][8] ), .S0(n5812), .S1(n5906), .Q(n4753) );
  MUX41X1 U5712 ( .IN1(\FIFO[0][8] ), .IN3(\FIFO[2][8] ), .IN2(\FIFO[1][8] ), 
        .IN4(\FIFO[3][8] ), .S0(n5812), .S1(n5906), .Q(n4754) );
  MUX41X1 U5713 ( .IN1(n4754), .IN3(n4752), .IN2(n4753), .IN4(n4751), .S0(
        n5740), .S1(n5778), .Q(n4755) );
  MUX41X1 U5714 ( .IN1(n4755), .IN3(n4745), .IN2(n4750), .IN4(n4740), .S0(
        n5727), .S1(n5731), .Q(n4756) );
  MUX21X1 U5715 ( .IN1(n4756), .IN2(n4735), .S(n5723), .Q(N242) );
  MUX41X1 U5716 ( .IN1(\FIFO[124][9] ), .IN3(\FIFO[126][9] ), .IN2(
        \FIFO[125][9] ), .IN4(\FIFO[127][9] ), .S0(n5812), .S1(n5906), .Q(
        n4757) );
  MUX41X1 U5717 ( .IN1(\FIFO[120][9] ), .IN3(\FIFO[122][9] ), .IN2(
        \FIFO[121][9] ), .IN4(\FIFO[123][9] ), .S0(n5812), .S1(n5906), .Q(
        n4758) );
  MUX41X1 U5718 ( .IN1(\FIFO[116][9] ), .IN3(\FIFO[118][9] ), .IN2(
        \FIFO[117][9] ), .IN4(\FIFO[119][9] ), .S0(n5812), .S1(n5906), .Q(
        n4759) );
  MUX41X1 U5719 ( .IN1(\FIFO[112][9] ), .IN3(\FIFO[114][9] ), .IN2(
        \FIFO[113][9] ), .IN4(\FIFO[115][9] ), .S0(n5812), .S1(n5906), .Q(
        n4760) );
  MUX41X1 U5720 ( .IN1(n4760), .IN3(n4758), .IN2(n4759), .IN4(n4757), .S0(
        n5740), .S1(n5778), .Q(n4761) );
  MUX41X1 U5721 ( .IN1(\FIFO[108][9] ), .IN3(\FIFO[110][9] ), .IN2(
        \FIFO[109][9] ), .IN4(\FIFO[111][9] ), .S0(n5813), .S1(n5907), .Q(
        n4762) );
  MUX41X1 U5722 ( .IN1(\FIFO[104][9] ), .IN3(\FIFO[106][9] ), .IN2(
        \FIFO[105][9] ), .IN4(\FIFO[107][9] ), .S0(n5813), .S1(n5907), .Q(
        n4763) );
  MUX41X1 U5723 ( .IN1(\FIFO[100][9] ), .IN3(\FIFO[102][9] ), .IN2(
        \FIFO[101][9] ), .IN4(\FIFO[103][9] ), .S0(n5813), .S1(n5907), .Q(
        n4764) );
  MUX41X1 U5724 ( .IN1(\FIFO[96][9] ), .IN3(\FIFO[98][9] ), .IN2(\FIFO[97][9] ), .IN4(\FIFO[99][9] ), .S0(n5813), .S1(n5907), .Q(n4765) );
  MUX41X1 U5725 ( .IN1(n4765), .IN3(n4763), .IN2(n4764), .IN4(n4762), .S0(
        n5740), .S1(n5781), .Q(n4766) );
  MUX41X1 U5726 ( .IN1(\FIFO[92][9] ), .IN3(\FIFO[94][9] ), .IN2(\FIFO[93][9] ), .IN4(\FIFO[95][9] ), .S0(n5813), .S1(n5907), .Q(n4767) );
  MUX41X1 U5727 ( .IN1(\FIFO[88][9] ), .IN3(\FIFO[90][9] ), .IN2(\FIFO[89][9] ), .IN4(\FIFO[91][9] ), .S0(n5813), .S1(n5907), .Q(n4768) );
  MUX41X1 U5728 ( .IN1(\FIFO[84][9] ), .IN3(\FIFO[86][9] ), .IN2(\FIFO[85][9] ), .IN4(\FIFO[87][9] ), .S0(n5813), .S1(n5907), .Q(n4769) );
  MUX41X1 U5729 ( .IN1(\FIFO[80][9] ), .IN3(\FIFO[82][9] ), .IN2(\FIFO[81][9] ), .IN4(\FIFO[83][9] ), .S0(n5813), .S1(n5907), .Q(n4770) );
  MUX41X1 U5730 ( .IN1(n4770), .IN3(n4768), .IN2(n4769), .IN4(n4767), .S0(
        n5740), .S1(n5776), .Q(n4771) );
  MUX41X1 U5731 ( .IN1(\FIFO[76][9] ), .IN3(\FIFO[78][9] ), .IN2(\FIFO[77][9] ), .IN4(\FIFO[79][9] ), .S0(n5813), .S1(n5907), .Q(n4772) );
  MUX41X1 U5732 ( .IN1(\FIFO[72][9] ), .IN3(\FIFO[74][9] ), .IN2(\FIFO[73][9] ), .IN4(\FIFO[75][9] ), .S0(n5813), .S1(n5907), .Q(n4773) );
  MUX41X1 U5733 ( .IN1(\FIFO[68][9] ), .IN3(\FIFO[70][9] ), .IN2(\FIFO[69][9] ), .IN4(\FIFO[71][9] ), .S0(n5813), .S1(n5907), .Q(n4774) );
  MUX41X1 U5734 ( .IN1(\FIFO[64][9] ), .IN3(\FIFO[66][9] ), .IN2(\FIFO[65][9] ), .IN4(\FIFO[67][9] ), .S0(n5813), .S1(n5907), .Q(n4775) );
  MUX41X1 U5735 ( .IN1(n4775), .IN3(n4773), .IN2(n4774), .IN4(n4772), .S0(
        n5740), .S1(n5779), .Q(n4776) );
  MUX41X1 U5736 ( .IN1(n4776), .IN3(n4766), .IN2(n4771), .IN4(n4761), .S0(
        n5727), .S1(n5731), .Q(n4777) );
  MUX41X1 U5737 ( .IN1(\FIFO[60][9] ), .IN3(\FIFO[62][9] ), .IN2(\FIFO[61][9] ), .IN4(\FIFO[63][9] ), .S0(n5814), .S1(n5908), .Q(n4778) );
  MUX41X1 U5738 ( .IN1(\FIFO[56][9] ), .IN3(\FIFO[58][9] ), .IN2(\FIFO[57][9] ), .IN4(\FIFO[59][9] ), .S0(n5814), .S1(n5908), .Q(n4779) );
  MUX41X1 U5739 ( .IN1(\FIFO[52][9] ), .IN3(\FIFO[54][9] ), .IN2(\FIFO[53][9] ), .IN4(\FIFO[55][9] ), .S0(n5814), .S1(n5908), .Q(n4780) );
  MUX41X1 U5740 ( .IN1(\FIFO[48][9] ), .IN3(\FIFO[50][9] ), .IN2(\FIFO[49][9] ), .IN4(\FIFO[51][9] ), .S0(n5814), .S1(n5908), .Q(n4781) );
  MUX41X1 U5741 ( .IN1(n4781), .IN3(n4779), .IN2(n4780), .IN4(n4778), .S0(
        n5741), .S1(n5760), .Q(n4782) );
  MUX41X1 U5742 ( .IN1(\FIFO[44][9] ), .IN3(\FIFO[46][9] ), .IN2(\FIFO[45][9] ), .IN4(\FIFO[47][9] ), .S0(n5814), .S1(n5908), .Q(n4783) );
  MUX41X1 U5743 ( .IN1(\FIFO[40][9] ), .IN3(\FIFO[42][9] ), .IN2(\FIFO[41][9] ), .IN4(\FIFO[43][9] ), .S0(n5814), .S1(n5908), .Q(n4784) );
  MUX41X1 U5744 ( .IN1(\FIFO[36][9] ), .IN3(\FIFO[38][9] ), .IN2(\FIFO[37][9] ), .IN4(\FIFO[39][9] ), .S0(n5814), .S1(n5908), .Q(n4785) );
  MUX41X1 U5745 ( .IN1(\FIFO[32][9] ), .IN3(\FIFO[34][9] ), .IN2(\FIFO[33][9] ), .IN4(\FIFO[35][9] ), .S0(n5814), .S1(n5908), .Q(n4786) );
  MUX41X1 U5746 ( .IN1(n4786), .IN3(n4784), .IN2(n4785), .IN4(n4783), .S0(
        n5741), .S1(n5760), .Q(n4787) );
  MUX41X1 U5747 ( .IN1(\FIFO[28][9] ), .IN3(\FIFO[30][9] ), .IN2(\FIFO[29][9] ), .IN4(\FIFO[31][9] ), .S0(n5814), .S1(n5908), .Q(n4788) );
  MUX41X1 U5748 ( .IN1(\FIFO[24][9] ), .IN3(\FIFO[26][9] ), .IN2(\FIFO[25][9] ), .IN4(\FIFO[27][9] ), .S0(n5814), .S1(n5908), .Q(n4789) );
  MUX41X1 U5749 ( .IN1(\FIFO[20][9] ), .IN3(\FIFO[22][9] ), .IN2(\FIFO[21][9] ), .IN4(\FIFO[23][9] ), .S0(n5814), .S1(n5908), .Q(n4790) );
  MUX41X1 U5750 ( .IN1(\FIFO[16][9] ), .IN3(\FIFO[18][9] ), .IN2(\FIFO[17][9] ), .IN4(\FIFO[19][9] ), .S0(n5814), .S1(n5908), .Q(n4791) );
  MUX41X1 U5751 ( .IN1(n4791), .IN3(n4789), .IN2(n4790), .IN4(n4788), .S0(
        n5741), .S1(n5760), .Q(n4792) );
  MUX41X1 U5752 ( .IN1(\FIFO[12][9] ), .IN3(\FIFO[14][9] ), .IN2(\FIFO[13][9] ), .IN4(\FIFO[15][9] ), .S0(n5815), .S1(n5909), .Q(n4793) );
  MUX41X1 U5753 ( .IN1(\FIFO[8][9] ), .IN3(\FIFO[10][9] ), .IN2(\FIFO[9][9] ), 
        .IN4(\FIFO[11][9] ), .S0(n5815), .S1(n5909), .Q(n4794) );
  MUX41X1 U5754 ( .IN1(\FIFO[4][9] ), .IN3(\FIFO[6][9] ), .IN2(\FIFO[5][9] ), 
        .IN4(\FIFO[7][9] ), .S0(n5815), .S1(n5909), .Q(n4795) );
  MUX41X1 U5755 ( .IN1(\FIFO[0][9] ), .IN3(\FIFO[2][9] ), .IN2(\FIFO[1][9] ), 
        .IN4(\FIFO[3][9] ), .S0(n5815), .S1(n5909), .Q(n4796) );
  MUX41X1 U5756 ( .IN1(n4796), .IN3(n4794), .IN2(n4795), .IN4(n4793), .S0(
        n5741), .S1(n5760), .Q(n4797) );
  MUX41X1 U5757 ( .IN1(n4797), .IN3(n4787), .IN2(n4792), .IN4(n4782), .S0(
        n5727), .S1(n5731), .Q(n4798) );
  MUX21X1 U5758 ( .IN1(n4798), .IN2(n4777), .S(n5723), .Q(N241) );
  MUX41X1 U5759 ( .IN1(\FIFO[124][10] ), .IN3(\FIFO[126][10] ), .IN2(
        \FIFO[125][10] ), .IN4(\FIFO[127][10] ), .S0(n5815), .S1(n5909), .Q(
        n4799) );
  MUX41X1 U5760 ( .IN1(\FIFO[120][10] ), .IN3(\FIFO[122][10] ), .IN2(
        \FIFO[121][10] ), .IN4(\FIFO[123][10] ), .S0(n5815), .S1(n5909), .Q(
        n4800) );
  MUX41X1 U5761 ( .IN1(\FIFO[116][10] ), .IN3(\FIFO[118][10] ), .IN2(
        \FIFO[117][10] ), .IN4(\FIFO[119][10] ), .S0(n5815), .S1(n5909), .Q(
        n4801) );
  MUX41X1 U5762 ( .IN1(\FIFO[112][10] ), .IN3(\FIFO[114][10] ), .IN2(
        \FIFO[113][10] ), .IN4(\FIFO[115][10] ), .S0(n5815), .S1(n5909), .Q(
        n4802) );
  MUX41X1 U5763 ( .IN1(n4802), .IN3(n4800), .IN2(n4801), .IN4(n4799), .S0(
        n5741), .S1(n5760), .Q(n4803) );
  MUX41X1 U5764 ( .IN1(\FIFO[108][10] ), .IN3(\FIFO[110][10] ), .IN2(
        \FIFO[109][10] ), .IN4(\FIFO[111][10] ), .S0(n5815), .S1(n5909), .Q(
        n4804) );
  MUX41X1 U5765 ( .IN1(\FIFO[104][10] ), .IN3(\FIFO[106][10] ), .IN2(
        \FIFO[105][10] ), .IN4(\FIFO[107][10] ), .S0(n5815), .S1(n5909), .Q(
        n4805) );
  MUX41X1 U5766 ( .IN1(\FIFO[100][10] ), .IN3(\FIFO[102][10] ), .IN2(
        \FIFO[101][10] ), .IN4(\FIFO[103][10] ), .S0(n5815), .S1(n5909), .Q(
        n4806) );
  MUX41X1 U5767 ( .IN1(\FIFO[96][10] ), .IN3(\FIFO[98][10] ), .IN2(
        \FIFO[97][10] ), .IN4(\FIFO[99][10] ), .S0(n5815), .S1(n5909), .Q(
        n4807) );
  MUX41X1 U5768 ( .IN1(n4807), .IN3(n4805), .IN2(n4806), .IN4(n4804), .S0(
        n5741), .S1(n5760), .Q(n4808) );
  MUX41X1 U5769 ( .IN1(\FIFO[92][10] ), .IN3(\FIFO[94][10] ), .IN2(
        \FIFO[93][10] ), .IN4(\FIFO[95][10] ), .S0(n5816), .S1(n5910), .Q(
        n4809) );
  MUX41X1 U5770 ( .IN1(\FIFO[88][10] ), .IN3(\FIFO[90][10] ), .IN2(
        \FIFO[89][10] ), .IN4(\FIFO[91][10] ), .S0(n5816), .S1(n5910), .Q(
        n4810) );
  MUX41X1 U5771 ( .IN1(\FIFO[84][10] ), .IN3(\FIFO[86][10] ), .IN2(
        \FIFO[85][10] ), .IN4(\FIFO[87][10] ), .S0(n5816), .S1(n5910), .Q(
        n4811) );
  MUX41X1 U5772 ( .IN1(\FIFO[80][10] ), .IN3(\FIFO[82][10] ), .IN2(
        \FIFO[81][10] ), .IN4(\FIFO[83][10] ), .S0(n5816), .S1(n5910), .Q(
        n4812) );
  MUX41X1 U5773 ( .IN1(n4812), .IN3(n4810), .IN2(n4811), .IN4(n4809), .S0(
        n5741), .S1(n5760), .Q(n4813) );
  MUX41X1 U5774 ( .IN1(\FIFO[76][10] ), .IN3(\FIFO[78][10] ), .IN2(
        \FIFO[77][10] ), .IN4(\FIFO[79][10] ), .S0(n5816), .S1(n5910), .Q(
        n4814) );
  MUX41X1 U5775 ( .IN1(\FIFO[72][10] ), .IN3(\FIFO[74][10] ), .IN2(
        \FIFO[73][10] ), .IN4(\FIFO[75][10] ), .S0(n5816), .S1(n5910), .Q(
        n4815) );
  MUX41X1 U5776 ( .IN1(\FIFO[68][10] ), .IN3(\FIFO[70][10] ), .IN2(
        \FIFO[69][10] ), .IN4(\FIFO[71][10] ), .S0(n5816), .S1(n5910), .Q(
        n4816) );
  MUX41X1 U5777 ( .IN1(\FIFO[64][10] ), .IN3(\FIFO[66][10] ), .IN2(
        \FIFO[65][10] ), .IN4(\FIFO[67][10] ), .S0(n5816), .S1(n5910), .Q(
        n4817) );
  MUX41X1 U5778 ( .IN1(n4817), .IN3(n4815), .IN2(n4816), .IN4(n4814), .S0(
        n5741), .S1(n5760), .Q(n4818) );
  MUX41X1 U5779 ( .IN1(n4818), .IN3(n4808), .IN2(n4813), .IN4(n4803), .S0(
        n5727), .S1(n5731), .Q(n4819) );
  MUX41X1 U5780 ( .IN1(\FIFO[60][10] ), .IN3(\FIFO[62][10] ), .IN2(
        \FIFO[61][10] ), .IN4(\FIFO[63][10] ), .S0(n5816), .S1(n5910), .Q(
        n4820) );
  MUX41X1 U5781 ( .IN1(\FIFO[56][10] ), .IN3(\FIFO[58][10] ), .IN2(
        \FIFO[57][10] ), .IN4(\FIFO[59][10] ), .S0(n5816), .S1(n5910), .Q(
        n4821) );
  MUX41X1 U5782 ( .IN1(\FIFO[52][10] ), .IN3(\FIFO[54][10] ), .IN2(
        \FIFO[53][10] ), .IN4(\FIFO[55][10] ), .S0(n5816), .S1(n5910), .Q(
        n4822) );
  MUX41X1 U5783 ( .IN1(\FIFO[48][10] ), .IN3(\FIFO[50][10] ), .IN2(
        \FIFO[49][10] ), .IN4(\FIFO[51][10] ), .S0(n5816), .S1(n5910), .Q(
        n4823) );
  MUX41X1 U5784 ( .IN1(n4823), .IN3(n4821), .IN2(n4822), .IN4(n4820), .S0(
        n5741), .S1(n5760), .Q(n4824) );
  MUX41X1 U5785 ( .IN1(\FIFO[44][10] ), .IN3(\FIFO[46][10] ), .IN2(
        \FIFO[45][10] ), .IN4(\FIFO[47][10] ), .S0(n5817), .S1(n5911), .Q(
        n4825) );
  MUX41X1 U5786 ( .IN1(\FIFO[40][10] ), .IN3(\FIFO[42][10] ), .IN2(
        \FIFO[41][10] ), .IN4(\FIFO[43][10] ), .S0(n5817), .S1(n5911), .Q(
        n4826) );
  MUX41X1 U5787 ( .IN1(\FIFO[36][10] ), .IN3(\FIFO[38][10] ), .IN2(
        \FIFO[37][10] ), .IN4(\FIFO[39][10] ), .S0(n5817), .S1(n5911), .Q(
        n4827) );
  MUX41X1 U5788 ( .IN1(\FIFO[32][10] ), .IN3(\FIFO[34][10] ), .IN2(
        \FIFO[33][10] ), .IN4(\FIFO[35][10] ), .S0(n5817), .S1(n5911), .Q(
        n4828) );
  MUX41X1 U5789 ( .IN1(n4828), .IN3(n4826), .IN2(n4827), .IN4(n4825), .S0(
        n5741), .S1(n5760), .Q(n4829) );
  MUX41X1 U5790 ( .IN1(\FIFO[28][10] ), .IN3(\FIFO[30][10] ), .IN2(
        \FIFO[29][10] ), .IN4(\FIFO[31][10] ), .S0(n5817), .S1(n5911), .Q(
        n4830) );
  MUX41X1 U5791 ( .IN1(\FIFO[24][10] ), .IN3(\FIFO[26][10] ), .IN2(
        \FIFO[25][10] ), .IN4(\FIFO[27][10] ), .S0(n5817), .S1(n5911), .Q(
        n4831) );
  MUX41X1 U5792 ( .IN1(\FIFO[20][10] ), .IN3(\FIFO[22][10] ), .IN2(
        \FIFO[21][10] ), .IN4(\FIFO[23][10] ), .S0(n5817), .S1(n5911), .Q(
        n4832) );
  MUX41X1 U5793 ( .IN1(\FIFO[16][10] ), .IN3(\FIFO[18][10] ), .IN2(
        \FIFO[17][10] ), .IN4(\FIFO[19][10] ), .S0(n5817), .S1(n5911), .Q(
        n4833) );
  MUX41X1 U5794 ( .IN1(n4833), .IN3(n4831), .IN2(n4832), .IN4(n4830), .S0(
        n5741), .S1(n5760), .Q(n4834) );
  MUX41X1 U5795 ( .IN1(\FIFO[12][10] ), .IN3(\FIFO[14][10] ), .IN2(
        \FIFO[13][10] ), .IN4(\FIFO[15][10] ), .S0(n5817), .S1(n5911), .Q(
        n4835) );
  MUX41X1 U5796 ( .IN1(\FIFO[8][10] ), .IN3(\FIFO[10][10] ), .IN2(
        \FIFO[9][10] ), .IN4(\FIFO[11][10] ), .S0(n5817), .S1(n5911), .Q(n4836) );
  MUX41X1 U5797 ( .IN1(\FIFO[4][10] ), .IN3(\FIFO[6][10] ), .IN2(\FIFO[5][10] ), .IN4(\FIFO[7][10] ), .S0(n5817), .S1(n5911), .Q(n4837) );
  MUX41X1 U5798 ( .IN1(\FIFO[0][10] ), .IN3(\FIFO[2][10] ), .IN2(\FIFO[1][10] ), .IN4(\FIFO[3][10] ), .S0(n5817), .S1(n5911), .Q(n4838) );
  MUX41X1 U5799 ( .IN1(n4838), .IN3(n4836), .IN2(n4837), .IN4(n4835), .S0(
        n5741), .S1(n5760), .Q(n4839) );
  MUX41X1 U5800 ( .IN1(n4839), .IN3(n4829), .IN2(n4834), .IN4(n4824), .S0(
        n5727), .S1(n5731), .Q(n4840) );
  MUX21X1 U5801 ( .IN1(n4840), .IN2(n4819), .S(n5723), .Q(N240) );
  MUX41X1 U5802 ( .IN1(\FIFO[124][11] ), .IN3(\FIFO[126][11] ), .IN2(
        \FIFO[125][11] ), .IN4(\FIFO[127][11] ), .S0(n5818), .S1(n5912), .Q(
        n4841) );
  MUX41X1 U5803 ( .IN1(\FIFO[120][11] ), .IN3(\FIFO[122][11] ), .IN2(
        \FIFO[121][11] ), .IN4(\FIFO[123][11] ), .S0(n5818), .S1(n5912), .Q(
        n4842) );
  MUX41X1 U5804 ( .IN1(\FIFO[116][11] ), .IN3(\FIFO[118][11] ), .IN2(
        \FIFO[117][11] ), .IN4(\FIFO[119][11] ), .S0(n5818), .S1(n5912), .Q(
        n4843) );
  MUX41X1 U5805 ( .IN1(\FIFO[112][11] ), .IN3(\FIFO[114][11] ), .IN2(
        \FIFO[113][11] ), .IN4(\FIFO[115][11] ), .S0(n5818), .S1(n5912), .Q(
        n4844) );
  MUX41X1 U5806 ( .IN1(n4844), .IN3(n4842), .IN2(n4843), .IN4(n4841), .S0(
        n5742), .S1(n5761), .Q(n4845) );
  MUX41X1 U5807 ( .IN1(\FIFO[108][11] ), .IN3(\FIFO[110][11] ), .IN2(
        \FIFO[109][11] ), .IN4(\FIFO[111][11] ), .S0(n5818), .S1(n5912), .Q(
        n4846) );
  MUX41X1 U5808 ( .IN1(\FIFO[104][11] ), .IN3(\FIFO[106][11] ), .IN2(
        \FIFO[105][11] ), .IN4(\FIFO[107][11] ), .S0(n5818), .S1(n5912), .Q(
        n4847) );
  MUX41X1 U5809 ( .IN1(\FIFO[100][11] ), .IN3(\FIFO[102][11] ), .IN2(
        \FIFO[101][11] ), .IN4(\FIFO[103][11] ), .S0(n5818), .S1(n5912), .Q(
        n4848) );
  MUX41X1 U5810 ( .IN1(\FIFO[96][11] ), .IN3(\FIFO[98][11] ), .IN2(
        \FIFO[97][11] ), .IN4(\FIFO[99][11] ), .S0(n5818), .S1(n5912), .Q(
        n4849) );
  MUX41X1 U5811 ( .IN1(n4849), .IN3(n4847), .IN2(n4848), .IN4(n4846), .S0(
        n5742), .S1(n5761), .Q(n4850) );
  MUX41X1 U5812 ( .IN1(\FIFO[92][11] ), .IN3(\FIFO[94][11] ), .IN2(
        \FIFO[93][11] ), .IN4(\FIFO[95][11] ), .S0(n5818), .S1(n5912), .Q(
        n4851) );
  MUX41X1 U5813 ( .IN1(\FIFO[88][11] ), .IN3(\FIFO[90][11] ), .IN2(
        \FIFO[89][11] ), .IN4(\FIFO[91][11] ), .S0(n5818), .S1(n5912), .Q(
        n4852) );
  MUX41X1 U5814 ( .IN1(\FIFO[84][11] ), .IN3(\FIFO[86][11] ), .IN2(
        \FIFO[85][11] ), .IN4(\FIFO[87][11] ), .S0(n5818), .S1(n5912), .Q(
        n4853) );
  MUX41X1 U5815 ( .IN1(\FIFO[80][11] ), .IN3(\FIFO[82][11] ), .IN2(
        \FIFO[81][11] ), .IN4(\FIFO[83][11] ), .S0(n5818), .S1(n5912), .Q(
        n4854) );
  MUX41X1 U5816 ( .IN1(n4854), .IN3(n4852), .IN2(n4853), .IN4(n4851), .S0(
        n5742), .S1(n5761), .Q(n4855) );
  MUX41X1 U5817 ( .IN1(\FIFO[76][11] ), .IN3(\FIFO[78][11] ), .IN2(
        \FIFO[77][11] ), .IN4(\FIFO[79][11] ), .S0(n5819), .S1(n5913), .Q(
        n4856) );
  MUX41X1 U5818 ( .IN1(\FIFO[72][11] ), .IN3(\FIFO[74][11] ), .IN2(
        \FIFO[73][11] ), .IN4(\FIFO[75][11] ), .S0(n5819), .S1(n5913), .Q(
        n4857) );
  MUX41X1 U5819 ( .IN1(\FIFO[68][11] ), .IN3(\FIFO[70][11] ), .IN2(
        \FIFO[69][11] ), .IN4(\FIFO[71][11] ), .S0(n5819), .S1(n5913), .Q(
        n4858) );
  MUX41X1 U5820 ( .IN1(\FIFO[64][11] ), .IN3(\FIFO[66][11] ), .IN2(
        \FIFO[65][11] ), .IN4(\FIFO[67][11] ), .S0(n5819), .S1(n5913), .Q(
        n4859) );
  MUX41X1 U5821 ( .IN1(n4859), .IN3(n4857), .IN2(n4858), .IN4(n4856), .S0(
        n5742), .S1(n5761), .Q(n4860) );
  MUX41X1 U5822 ( .IN1(n4860), .IN3(n4850), .IN2(n4855), .IN4(n4845), .S0(
        n5727), .S1(n5731), .Q(n4861) );
  MUX41X1 U5823 ( .IN1(\FIFO[60][11] ), .IN3(\FIFO[62][11] ), .IN2(
        \FIFO[61][11] ), .IN4(\FIFO[63][11] ), .S0(n5819), .S1(n5913), .Q(
        n4862) );
  MUX41X1 U5824 ( .IN1(\FIFO[56][11] ), .IN3(\FIFO[58][11] ), .IN2(
        \FIFO[57][11] ), .IN4(\FIFO[59][11] ), .S0(n5819), .S1(n5913), .Q(
        n4863) );
  MUX41X1 U5825 ( .IN1(\FIFO[52][11] ), .IN3(\FIFO[54][11] ), .IN2(
        \FIFO[53][11] ), .IN4(\FIFO[55][11] ), .S0(n5819), .S1(n5913), .Q(
        n4864) );
  MUX41X1 U5826 ( .IN1(\FIFO[48][11] ), .IN3(\FIFO[50][11] ), .IN2(
        \FIFO[49][11] ), .IN4(\FIFO[51][11] ), .S0(n5819), .S1(n5913), .Q(
        n4865) );
  MUX41X1 U5827 ( .IN1(n4865), .IN3(n4863), .IN2(n4864), .IN4(n4862), .S0(
        n5742), .S1(n5761), .Q(n4866) );
  MUX41X1 U5828 ( .IN1(\FIFO[44][11] ), .IN3(\FIFO[46][11] ), .IN2(
        \FIFO[45][11] ), .IN4(\FIFO[47][11] ), .S0(n5819), .S1(n5913), .Q(
        n4867) );
  MUX41X1 U5829 ( .IN1(\FIFO[40][11] ), .IN3(\FIFO[42][11] ), .IN2(
        \FIFO[41][11] ), .IN4(\FIFO[43][11] ), .S0(n5819), .S1(n5913), .Q(
        n4868) );
  MUX41X1 U5830 ( .IN1(\FIFO[36][11] ), .IN3(\FIFO[38][11] ), .IN2(
        \FIFO[37][11] ), .IN4(\FIFO[39][11] ), .S0(n5819), .S1(n5913), .Q(
        n4869) );
  MUX41X1 U5831 ( .IN1(\FIFO[32][11] ), .IN3(\FIFO[34][11] ), .IN2(
        \FIFO[33][11] ), .IN4(\FIFO[35][11] ), .S0(n5819), .S1(n5913), .Q(
        n4870) );
  MUX41X1 U5832 ( .IN1(n4870), .IN3(n4868), .IN2(n4869), .IN4(n4867), .S0(
        n5742), .S1(n5761), .Q(n4871) );
  MUX41X1 U5833 ( .IN1(\FIFO[28][11] ), .IN3(\FIFO[30][11] ), .IN2(
        \FIFO[29][11] ), .IN4(\FIFO[31][11] ), .S0(n5820), .S1(n5914), .Q(
        n4872) );
  MUX41X1 U5834 ( .IN1(\FIFO[24][11] ), .IN3(\FIFO[26][11] ), .IN2(
        \FIFO[25][11] ), .IN4(\FIFO[27][11] ), .S0(n5820), .S1(n5914), .Q(
        n4873) );
  MUX41X1 U5835 ( .IN1(\FIFO[20][11] ), .IN3(\FIFO[22][11] ), .IN2(
        \FIFO[21][11] ), .IN4(\FIFO[23][11] ), .S0(n5820), .S1(n5914), .Q(
        n4874) );
  MUX41X1 U5836 ( .IN1(\FIFO[16][11] ), .IN3(\FIFO[18][11] ), .IN2(
        \FIFO[17][11] ), .IN4(\FIFO[19][11] ), .S0(n5820), .S1(n5914), .Q(
        n4875) );
  MUX41X1 U5837 ( .IN1(n4875), .IN3(n4873), .IN2(n4874), .IN4(n4872), .S0(
        n5742), .S1(n5761), .Q(n4876) );
  MUX41X1 U5838 ( .IN1(\FIFO[12][11] ), .IN3(\FIFO[14][11] ), .IN2(
        \FIFO[13][11] ), .IN4(\FIFO[15][11] ), .S0(n5820), .S1(n5914), .Q(
        n4877) );
  MUX41X1 U5839 ( .IN1(\FIFO[8][11] ), .IN3(\FIFO[10][11] ), .IN2(
        \FIFO[9][11] ), .IN4(\FIFO[11][11] ), .S0(n5820), .S1(n5914), .Q(n4878) );
  MUX41X1 U5840 ( .IN1(\FIFO[4][11] ), .IN3(\FIFO[6][11] ), .IN2(\FIFO[5][11] ), .IN4(\FIFO[7][11] ), .S0(n5820), .S1(n5914), .Q(n4879) );
  MUX41X1 U5841 ( .IN1(\FIFO[0][11] ), .IN3(\FIFO[2][11] ), .IN2(\FIFO[1][11] ), .IN4(\FIFO[3][11] ), .S0(n5820), .S1(n5914), .Q(n4880) );
  MUX41X1 U5842 ( .IN1(n4880), .IN3(n4878), .IN2(n4879), .IN4(n4877), .S0(
        n5742), .S1(n5761), .Q(n4881) );
  MUX41X1 U5843 ( .IN1(n4881), .IN3(n4871), .IN2(n4876), .IN4(n4866), .S0(
        n5727), .S1(n5731), .Q(n4882) );
  MUX21X1 U5844 ( .IN1(n4882), .IN2(n4861), .S(n5723), .Q(N239) );
  MUX41X1 U5845 ( .IN1(\FIFO[124][12] ), .IN3(\FIFO[126][12] ), .IN2(
        \FIFO[125][12] ), .IN4(\FIFO[127][12] ), .S0(n5820), .S1(n5914), .Q(
        n4883) );
  MUX41X1 U5846 ( .IN1(\FIFO[120][12] ), .IN3(\FIFO[122][12] ), .IN2(
        \FIFO[121][12] ), .IN4(\FIFO[123][12] ), .S0(n5820), .S1(n5914), .Q(
        n4884) );
  MUX41X1 U5847 ( .IN1(\FIFO[116][12] ), .IN3(\FIFO[118][12] ), .IN2(
        \FIFO[117][12] ), .IN4(\FIFO[119][12] ), .S0(n5820), .S1(n5914), .Q(
        n4885) );
  MUX41X1 U5848 ( .IN1(\FIFO[112][12] ), .IN3(\FIFO[114][12] ), .IN2(
        \FIFO[113][12] ), .IN4(\FIFO[115][12] ), .S0(n5820), .S1(n5914), .Q(
        n4886) );
  MUX41X1 U5849 ( .IN1(n4886), .IN3(n4884), .IN2(n4885), .IN4(n4883), .S0(
        n5742), .S1(n5761), .Q(n4887) );
  MUX41X1 U5850 ( .IN1(\FIFO[108][12] ), .IN3(\FIFO[110][12] ), .IN2(
        \FIFO[109][12] ), .IN4(\FIFO[111][12] ), .S0(n5821), .S1(n5915), .Q(
        n4888) );
  MUX41X1 U5851 ( .IN1(\FIFO[104][12] ), .IN3(\FIFO[106][12] ), .IN2(
        \FIFO[105][12] ), .IN4(\FIFO[107][12] ), .S0(n5821), .S1(n5915), .Q(
        n4889) );
  MUX41X1 U5852 ( .IN1(\FIFO[100][12] ), .IN3(\FIFO[102][12] ), .IN2(
        \FIFO[101][12] ), .IN4(\FIFO[103][12] ), .S0(n5821), .S1(n5915), .Q(
        n4890) );
  MUX41X1 U5853 ( .IN1(\FIFO[96][12] ), .IN3(\FIFO[98][12] ), .IN2(
        \FIFO[97][12] ), .IN4(\FIFO[99][12] ), .S0(n5821), .S1(n5915), .Q(
        n4891) );
  MUX41X1 U5854 ( .IN1(n4891), .IN3(n4889), .IN2(n4890), .IN4(n4888), .S0(
        n5742), .S1(n5761), .Q(n4892) );
  MUX41X1 U5855 ( .IN1(\FIFO[92][12] ), .IN3(\FIFO[94][12] ), .IN2(
        \FIFO[93][12] ), .IN4(\FIFO[95][12] ), .S0(n5821), .S1(n5915), .Q(
        n4893) );
  MUX41X1 U5856 ( .IN1(\FIFO[88][12] ), .IN3(\FIFO[90][12] ), .IN2(
        \FIFO[89][12] ), .IN4(\FIFO[91][12] ), .S0(n5821), .S1(n5915), .Q(
        n4894) );
  MUX41X1 U5857 ( .IN1(\FIFO[84][12] ), .IN3(\FIFO[86][12] ), .IN2(
        \FIFO[85][12] ), .IN4(\FIFO[87][12] ), .S0(n5821), .S1(n5915), .Q(
        n4895) );
  MUX41X1 U5858 ( .IN1(\FIFO[80][12] ), .IN3(\FIFO[82][12] ), .IN2(
        \FIFO[81][12] ), .IN4(\FIFO[83][12] ), .S0(n5821), .S1(n5915), .Q(
        n4896) );
  MUX41X1 U5859 ( .IN1(n4896), .IN3(n4894), .IN2(n4895), .IN4(n4893), .S0(
        n5742), .S1(n5761), .Q(n4897) );
  MUX41X1 U5860 ( .IN1(\FIFO[76][12] ), .IN3(\FIFO[78][12] ), .IN2(
        \FIFO[77][12] ), .IN4(\FIFO[79][12] ), .S0(n5821), .S1(n5915), .Q(
        n4898) );
  MUX41X1 U5861 ( .IN1(\FIFO[72][12] ), .IN3(\FIFO[74][12] ), .IN2(
        \FIFO[73][12] ), .IN4(\FIFO[75][12] ), .S0(n5821), .S1(n5915), .Q(
        n4899) );
  MUX41X1 U5862 ( .IN1(\FIFO[68][12] ), .IN3(\FIFO[70][12] ), .IN2(
        \FIFO[69][12] ), .IN4(\FIFO[71][12] ), .S0(n5821), .S1(n5915), .Q(
        n4900) );
  MUX41X1 U5863 ( .IN1(\FIFO[64][12] ), .IN3(\FIFO[66][12] ), .IN2(
        \FIFO[65][12] ), .IN4(\FIFO[67][12] ), .S0(n5821), .S1(n5915), .Q(
        n4901) );
  MUX41X1 U5864 ( .IN1(n4901), .IN3(n4899), .IN2(n4900), .IN4(n4898), .S0(
        n5742), .S1(n5761), .Q(n4902) );
  MUX41X1 U5865 ( .IN1(n4902), .IN3(n4892), .IN2(n4897), .IN4(n4887), .S0(
        n5727), .S1(n5731), .Q(n4903) );
  MUX41X1 U5866 ( .IN1(\FIFO[60][12] ), .IN3(\FIFO[62][12] ), .IN2(
        \FIFO[61][12] ), .IN4(\FIFO[63][12] ), .S0(n5822), .S1(n5916), .Q(
        n4904) );
  MUX41X1 U5867 ( .IN1(\FIFO[56][12] ), .IN3(\FIFO[58][12] ), .IN2(
        \FIFO[57][12] ), .IN4(\FIFO[59][12] ), .S0(n5822), .S1(n5916), .Q(
        n4905) );
  MUX41X1 U5868 ( .IN1(\FIFO[52][12] ), .IN3(\FIFO[54][12] ), .IN2(
        \FIFO[53][12] ), .IN4(\FIFO[55][12] ), .S0(n5822), .S1(n5916), .Q(
        n4906) );
  MUX41X1 U5869 ( .IN1(\FIFO[48][12] ), .IN3(\FIFO[50][12] ), .IN2(
        \FIFO[49][12] ), .IN4(\FIFO[51][12] ), .S0(n5822), .S1(n5916), .Q(
        n4907) );
  MUX41X1 U5870 ( .IN1(n4907), .IN3(n4905), .IN2(n4906), .IN4(n4904), .S0(
        n5743), .S1(n5762), .Q(n4908) );
  MUX41X1 U5871 ( .IN1(\FIFO[44][12] ), .IN3(\FIFO[46][12] ), .IN2(
        \FIFO[45][12] ), .IN4(\FIFO[47][12] ), .S0(n5822), .S1(n5916), .Q(
        n4909) );
  MUX41X1 U5872 ( .IN1(\FIFO[40][12] ), .IN3(\FIFO[42][12] ), .IN2(
        \FIFO[41][12] ), .IN4(\FIFO[43][12] ), .S0(n5822), .S1(n5916), .Q(
        n4910) );
  MUX41X1 U5873 ( .IN1(\FIFO[36][12] ), .IN3(\FIFO[38][12] ), .IN2(
        \FIFO[37][12] ), .IN4(\FIFO[39][12] ), .S0(n5822), .S1(n5916), .Q(
        n4911) );
  MUX41X1 U5874 ( .IN1(\FIFO[32][12] ), .IN3(\FIFO[34][12] ), .IN2(
        \FIFO[33][12] ), .IN4(\FIFO[35][12] ), .S0(n5822), .S1(n5916), .Q(
        n4912) );
  MUX41X1 U5875 ( .IN1(n4912), .IN3(n4910), .IN2(n4911), .IN4(n4909), .S0(
        n5743), .S1(n5762), .Q(n4913) );
  MUX41X1 U5876 ( .IN1(\FIFO[28][12] ), .IN3(\FIFO[30][12] ), .IN2(
        \FIFO[29][12] ), .IN4(\FIFO[31][12] ), .S0(n5822), .S1(n5916), .Q(
        n4914) );
  MUX41X1 U5877 ( .IN1(\FIFO[24][12] ), .IN3(\FIFO[26][12] ), .IN2(
        \FIFO[25][12] ), .IN4(\FIFO[27][12] ), .S0(n5822), .S1(n5916), .Q(
        n4915) );
  MUX41X1 U5878 ( .IN1(\FIFO[20][12] ), .IN3(\FIFO[22][12] ), .IN2(
        \FIFO[21][12] ), .IN4(\FIFO[23][12] ), .S0(n5822), .S1(n5916), .Q(
        n4916) );
  MUX41X1 U5879 ( .IN1(\FIFO[16][12] ), .IN3(\FIFO[18][12] ), .IN2(
        \FIFO[17][12] ), .IN4(\FIFO[19][12] ), .S0(n5822), .S1(n5916), .Q(
        n4917) );
  MUX41X1 U5880 ( .IN1(n4917), .IN3(n4915), .IN2(n4916), .IN4(n4914), .S0(
        n5743), .S1(n5762), .Q(n4918) );
  MUX41X1 U5881 ( .IN1(\FIFO[12][12] ), .IN3(\FIFO[14][12] ), .IN2(
        \FIFO[13][12] ), .IN4(\FIFO[15][12] ), .S0(n5823), .S1(n5917), .Q(
        n4919) );
  MUX41X1 U5882 ( .IN1(\FIFO[8][12] ), .IN3(\FIFO[10][12] ), .IN2(
        \FIFO[9][12] ), .IN4(\FIFO[11][12] ), .S0(n5823), .S1(n5917), .Q(n4920) );
  MUX41X1 U5883 ( .IN1(\FIFO[4][12] ), .IN3(\FIFO[6][12] ), .IN2(\FIFO[5][12] ), .IN4(\FIFO[7][12] ), .S0(n5823), .S1(n5917), .Q(n4921) );
  MUX41X1 U5884 ( .IN1(\FIFO[0][12] ), .IN3(\FIFO[2][12] ), .IN2(\FIFO[1][12] ), .IN4(\FIFO[3][12] ), .S0(n5823), .S1(n5917), .Q(n4922) );
  MUX41X1 U5885 ( .IN1(n4922), .IN3(n4920), .IN2(n4921), .IN4(n4919), .S0(
        n5743), .S1(n5762), .Q(n4923) );
  MUX41X1 U5886 ( .IN1(n4923), .IN3(n4913), .IN2(n4918), .IN4(n4908), .S0(
        n5727), .S1(n5731), .Q(n4924) );
  MUX21X1 U5887 ( .IN1(n4924), .IN2(n4903), .S(n5723), .Q(N238) );
  MUX41X1 U5888 ( .IN1(\FIFO[124][13] ), .IN3(\FIFO[126][13] ), .IN2(
        \FIFO[125][13] ), .IN4(\FIFO[127][13] ), .S0(n5823), .S1(n5917), .Q(
        n4925) );
  MUX41X1 U5889 ( .IN1(\FIFO[120][13] ), .IN3(\FIFO[122][13] ), .IN2(
        \FIFO[121][13] ), .IN4(\FIFO[123][13] ), .S0(n5823), .S1(n5917), .Q(
        n4926) );
  MUX41X1 U5890 ( .IN1(\FIFO[116][13] ), .IN3(\FIFO[118][13] ), .IN2(
        \FIFO[117][13] ), .IN4(\FIFO[119][13] ), .S0(n5823), .S1(n5917), .Q(
        n4927) );
  MUX41X1 U5891 ( .IN1(\FIFO[112][13] ), .IN3(\FIFO[114][13] ), .IN2(
        \FIFO[113][13] ), .IN4(\FIFO[115][13] ), .S0(n5823), .S1(n5917), .Q(
        n4928) );
  MUX41X1 U5892 ( .IN1(n4928), .IN3(n4926), .IN2(n4927), .IN4(n4925), .S0(
        n5743), .S1(n5762), .Q(n4929) );
  MUX41X1 U5893 ( .IN1(\FIFO[108][13] ), .IN3(\FIFO[110][13] ), .IN2(
        \FIFO[109][13] ), .IN4(\FIFO[111][13] ), .S0(n5823), .S1(n5917), .Q(
        n4930) );
  MUX41X1 U5894 ( .IN1(\FIFO[104][13] ), .IN3(\FIFO[106][13] ), .IN2(
        \FIFO[105][13] ), .IN4(\FIFO[107][13] ), .S0(n5823), .S1(n5917), .Q(
        n4931) );
  MUX41X1 U5895 ( .IN1(\FIFO[100][13] ), .IN3(\FIFO[102][13] ), .IN2(
        \FIFO[101][13] ), .IN4(\FIFO[103][13] ), .S0(n5823), .S1(n5917), .Q(
        n4932) );
  MUX41X1 U5896 ( .IN1(\FIFO[96][13] ), .IN3(\FIFO[98][13] ), .IN2(
        \FIFO[97][13] ), .IN4(\FIFO[99][13] ), .S0(n5823), .S1(n5917), .Q(
        n4933) );
  MUX41X1 U5897 ( .IN1(n4933), .IN3(n4931), .IN2(n4932), .IN4(n4930), .S0(
        n5743), .S1(n5762), .Q(n4934) );
  MUX41X1 U5898 ( .IN1(\FIFO[92][13] ), .IN3(\FIFO[94][13] ), .IN2(
        \FIFO[93][13] ), .IN4(\FIFO[95][13] ), .S0(n5824), .S1(n5918), .Q(
        n4935) );
  MUX41X1 U5899 ( .IN1(\FIFO[88][13] ), .IN3(\FIFO[90][13] ), .IN2(
        \FIFO[89][13] ), .IN4(\FIFO[91][13] ), .S0(n5824), .S1(n5918), .Q(
        n4936) );
  MUX41X1 U5900 ( .IN1(\FIFO[84][13] ), .IN3(\FIFO[86][13] ), .IN2(
        \FIFO[85][13] ), .IN4(\FIFO[87][13] ), .S0(n5824), .S1(n5918), .Q(
        n4937) );
  MUX41X1 U5901 ( .IN1(\FIFO[80][13] ), .IN3(\FIFO[82][13] ), .IN2(
        \FIFO[81][13] ), .IN4(\FIFO[83][13] ), .S0(n5824), .S1(n5918), .Q(
        n4938) );
  MUX41X1 U5902 ( .IN1(n4938), .IN3(n4936), .IN2(n4937), .IN4(n4935), .S0(
        n5743), .S1(n5762), .Q(n4939) );
  MUX41X1 U5903 ( .IN1(\FIFO[76][13] ), .IN3(\FIFO[78][13] ), .IN2(
        \FIFO[77][13] ), .IN4(\FIFO[79][13] ), .S0(n5824), .S1(n5918), .Q(
        n4940) );
  MUX41X1 U5904 ( .IN1(\FIFO[72][13] ), .IN3(\FIFO[74][13] ), .IN2(
        \FIFO[73][13] ), .IN4(\FIFO[75][13] ), .S0(n5824), .S1(n5918), .Q(
        n4941) );
  MUX41X1 U5905 ( .IN1(\FIFO[68][13] ), .IN3(\FIFO[70][13] ), .IN2(
        \FIFO[69][13] ), .IN4(\FIFO[71][13] ), .S0(n5824), .S1(n5918), .Q(
        n4942) );
  MUX41X1 U5906 ( .IN1(\FIFO[64][13] ), .IN3(\FIFO[66][13] ), .IN2(
        \FIFO[65][13] ), .IN4(\FIFO[67][13] ), .S0(n5824), .S1(n5918), .Q(
        n4943) );
  MUX41X1 U5907 ( .IN1(n4943), .IN3(n4941), .IN2(n4942), .IN4(n4940), .S0(
        n5743), .S1(n5762), .Q(n4944) );
  MUX41X1 U5908 ( .IN1(n4944), .IN3(n4934), .IN2(n4939), .IN4(n4929), .S0(
        n5727), .S1(n5731), .Q(n4945) );
  MUX41X1 U5909 ( .IN1(\FIFO[60][13] ), .IN3(\FIFO[62][13] ), .IN2(
        \FIFO[61][13] ), .IN4(\FIFO[63][13] ), .S0(n5824), .S1(n5918), .Q(
        n4946) );
  MUX41X1 U5910 ( .IN1(\FIFO[56][13] ), .IN3(\FIFO[58][13] ), .IN2(
        \FIFO[57][13] ), .IN4(\FIFO[59][13] ), .S0(n5824), .S1(n5918), .Q(
        n4947) );
  MUX41X1 U5911 ( .IN1(\FIFO[52][13] ), .IN3(\FIFO[54][13] ), .IN2(
        \FIFO[53][13] ), .IN4(\FIFO[55][13] ), .S0(n5824), .S1(n5918), .Q(
        n4948) );
  MUX41X1 U5912 ( .IN1(\FIFO[48][13] ), .IN3(\FIFO[50][13] ), .IN2(
        \FIFO[49][13] ), .IN4(\FIFO[51][13] ), .S0(n5824), .S1(n5918), .Q(
        n4949) );
  MUX41X1 U5913 ( .IN1(n4949), .IN3(n4947), .IN2(n4948), .IN4(n4946), .S0(
        n5743), .S1(n5762), .Q(n4950) );
  MUX41X1 U5914 ( .IN1(\FIFO[44][13] ), .IN3(\FIFO[46][13] ), .IN2(
        \FIFO[45][13] ), .IN4(\FIFO[47][13] ), .S0(n5825), .S1(n5919), .Q(
        n4951) );
  MUX41X1 U5915 ( .IN1(\FIFO[40][13] ), .IN3(\FIFO[42][13] ), .IN2(
        \FIFO[41][13] ), .IN4(\FIFO[43][13] ), .S0(n5825), .S1(n5919), .Q(
        n4952) );
  MUX41X1 U5916 ( .IN1(\FIFO[36][13] ), .IN3(\FIFO[38][13] ), .IN2(
        \FIFO[37][13] ), .IN4(\FIFO[39][13] ), .S0(n5825), .S1(n5919), .Q(
        n4953) );
  MUX41X1 U5917 ( .IN1(\FIFO[32][13] ), .IN3(\FIFO[34][13] ), .IN2(
        \FIFO[33][13] ), .IN4(\FIFO[35][13] ), .S0(n5825), .S1(n5919), .Q(
        n4954) );
  MUX41X1 U5918 ( .IN1(n4954), .IN3(n4952), .IN2(n4953), .IN4(n4951), .S0(
        n5743), .S1(n5762), .Q(n4955) );
  MUX41X1 U5919 ( .IN1(\FIFO[28][13] ), .IN3(\FIFO[30][13] ), .IN2(
        \FIFO[29][13] ), .IN4(\FIFO[31][13] ), .S0(n5825), .S1(n5919), .Q(
        n4956) );
  MUX41X1 U5920 ( .IN1(\FIFO[24][13] ), .IN3(\FIFO[26][13] ), .IN2(
        \FIFO[25][13] ), .IN4(\FIFO[27][13] ), .S0(n5825), .S1(n5919), .Q(
        n4957) );
  MUX41X1 U5921 ( .IN1(\FIFO[20][13] ), .IN3(\FIFO[22][13] ), .IN2(
        \FIFO[21][13] ), .IN4(\FIFO[23][13] ), .S0(n5825), .S1(n5919), .Q(
        n4958) );
  MUX41X1 U5922 ( .IN1(\FIFO[16][13] ), .IN3(\FIFO[18][13] ), .IN2(
        \FIFO[17][13] ), .IN4(\FIFO[19][13] ), .S0(n5825), .S1(n5919), .Q(
        n4959) );
  MUX41X1 U5923 ( .IN1(n4959), .IN3(n4957), .IN2(n4958), .IN4(n4956), .S0(
        n5743), .S1(n5762), .Q(n4960) );
  MUX41X1 U5924 ( .IN1(\FIFO[12][13] ), .IN3(\FIFO[14][13] ), .IN2(
        \FIFO[13][13] ), .IN4(\FIFO[15][13] ), .S0(n5825), .S1(n5919), .Q(
        n4961) );
  MUX41X1 U5925 ( .IN1(\FIFO[8][13] ), .IN3(\FIFO[10][13] ), .IN2(
        \FIFO[9][13] ), .IN4(\FIFO[11][13] ), .S0(n5825), .S1(n5919), .Q(n4962) );
  MUX41X1 U5926 ( .IN1(\FIFO[4][13] ), .IN3(\FIFO[6][13] ), .IN2(\FIFO[5][13] ), .IN4(\FIFO[7][13] ), .S0(n5825), .S1(n5919), .Q(n4963) );
  MUX41X1 U5927 ( .IN1(\FIFO[0][13] ), .IN3(\FIFO[2][13] ), .IN2(\FIFO[1][13] ), .IN4(\FIFO[3][13] ), .S0(n5825), .S1(n5919), .Q(n4964) );
  MUX41X1 U5928 ( .IN1(n4964), .IN3(n4962), .IN2(n4963), .IN4(n4961), .S0(
        n5743), .S1(n5762), .Q(n4965) );
  MUX41X1 U5929 ( .IN1(n4965), .IN3(n4955), .IN2(n4960), .IN4(n4950), .S0(
        n5727), .S1(n5731), .Q(n4966) );
  MUX21X1 U5930 ( .IN1(n4966), .IN2(n4945), .S(n5723), .Q(N237) );
  MUX41X1 U5931 ( .IN1(\FIFO[124][14] ), .IN3(\FIFO[126][14] ), .IN2(
        \FIFO[125][14] ), .IN4(\FIFO[127][14] ), .S0(n5826), .S1(n5920), .Q(
        n4967) );
  MUX41X1 U5932 ( .IN1(\FIFO[120][14] ), .IN3(\FIFO[122][14] ), .IN2(
        \FIFO[121][14] ), .IN4(\FIFO[123][14] ), .S0(n5826), .S1(n5920), .Q(
        n4968) );
  MUX41X1 U5933 ( .IN1(\FIFO[116][14] ), .IN3(\FIFO[118][14] ), .IN2(
        \FIFO[117][14] ), .IN4(\FIFO[119][14] ), .S0(n5826), .S1(n5920), .Q(
        n4969) );
  MUX41X1 U5934 ( .IN1(\FIFO[112][14] ), .IN3(\FIFO[114][14] ), .IN2(
        \FIFO[113][14] ), .IN4(\FIFO[115][14] ), .S0(n5826), .S1(n5920), .Q(
        n4970) );
  MUX41X1 U5935 ( .IN1(n4970), .IN3(n4968), .IN2(n4969), .IN4(n4967), .S0(
        n5744), .S1(n5763), .Q(n4971) );
  MUX41X1 U5936 ( .IN1(\FIFO[108][14] ), .IN3(\FIFO[110][14] ), .IN2(
        \FIFO[109][14] ), .IN4(\FIFO[111][14] ), .S0(n5826), .S1(n5920), .Q(
        n4972) );
  MUX41X1 U5937 ( .IN1(\FIFO[104][14] ), .IN3(\FIFO[106][14] ), .IN2(
        \FIFO[105][14] ), .IN4(\FIFO[107][14] ), .S0(n5826), .S1(n5920), .Q(
        n4973) );
  MUX41X1 U5938 ( .IN1(\FIFO[100][14] ), .IN3(\FIFO[102][14] ), .IN2(
        \FIFO[101][14] ), .IN4(\FIFO[103][14] ), .S0(n5826), .S1(n5920), .Q(
        n4974) );
  MUX41X1 U5939 ( .IN1(\FIFO[96][14] ), .IN3(\FIFO[98][14] ), .IN2(
        \FIFO[97][14] ), .IN4(\FIFO[99][14] ), .S0(n5826), .S1(n5920), .Q(
        n4975) );
  MUX41X1 U5940 ( .IN1(n4975), .IN3(n4973), .IN2(n4974), .IN4(n4972), .S0(
        n5744), .S1(n5763), .Q(n4976) );
  MUX41X1 U5941 ( .IN1(\FIFO[92][14] ), .IN3(\FIFO[94][14] ), .IN2(
        \FIFO[93][14] ), .IN4(\FIFO[95][14] ), .S0(n5826), .S1(n5920), .Q(
        n4977) );
  MUX41X1 U5942 ( .IN1(\FIFO[88][14] ), .IN3(\FIFO[90][14] ), .IN2(
        \FIFO[89][14] ), .IN4(\FIFO[91][14] ), .S0(n5826), .S1(n5920), .Q(
        n4978) );
  MUX41X1 U5943 ( .IN1(\FIFO[84][14] ), .IN3(\FIFO[86][14] ), .IN2(
        \FIFO[85][14] ), .IN4(\FIFO[87][14] ), .S0(n5826), .S1(n5920), .Q(
        n4979) );
  MUX41X1 U5944 ( .IN1(\FIFO[80][14] ), .IN3(\FIFO[82][14] ), .IN2(
        \FIFO[81][14] ), .IN4(\FIFO[83][14] ), .S0(n5826), .S1(n5920), .Q(
        n4980) );
  MUX41X1 U5945 ( .IN1(n4980), .IN3(n4978), .IN2(n4979), .IN4(n4977), .S0(
        n5744), .S1(n5763), .Q(n4981) );
  MUX41X1 U5946 ( .IN1(\FIFO[76][14] ), .IN3(\FIFO[78][14] ), .IN2(
        \FIFO[77][14] ), .IN4(\FIFO[79][14] ), .S0(n5827), .S1(n5921), .Q(
        n4982) );
  MUX41X1 U5947 ( .IN1(\FIFO[72][14] ), .IN3(\FIFO[74][14] ), .IN2(
        \FIFO[73][14] ), .IN4(\FIFO[75][14] ), .S0(n5827), .S1(n5921), .Q(
        n4983) );
  MUX41X1 U5948 ( .IN1(\FIFO[68][14] ), .IN3(\FIFO[70][14] ), .IN2(
        \FIFO[69][14] ), .IN4(\FIFO[71][14] ), .S0(n5827), .S1(n5921), .Q(
        n4984) );
  MUX41X1 U5949 ( .IN1(\FIFO[64][14] ), .IN3(\FIFO[66][14] ), .IN2(
        \FIFO[65][14] ), .IN4(\FIFO[67][14] ), .S0(n5827), .S1(n5921), .Q(
        n4985) );
  MUX41X1 U5950 ( .IN1(n4985), .IN3(n4983), .IN2(n4984), .IN4(n4982), .S0(
        n5744), .S1(n5763), .Q(n4986) );
  MUX41X1 U5951 ( .IN1(n4986), .IN3(n4976), .IN2(n4981), .IN4(n4971), .S0(
        n5728), .S1(n5732), .Q(n4987) );
  MUX41X1 U5952 ( .IN1(\FIFO[60][14] ), .IN3(\FIFO[62][14] ), .IN2(
        \FIFO[61][14] ), .IN4(\FIFO[63][14] ), .S0(n5827), .S1(n5921), .Q(
        n4988) );
  MUX41X1 U5953 ( .IN1(\FIFO[56][14] ), .IN3(\FIFO[58][14] ), .IN2(
        \FIFO[57][14] ), .IN4(\FIFO[59][14] ), .S0(n5827), .S1(n5921), .Q(
        n4989) );
  MUX41X1 U5954 ( .IN1(\FIFO[52][14] ), .IN3(\FIFO[54][14] ), .IN2(
        \FIFO[53][14] ), .IN4(\FIFO[55][14] ), .S0(n5827), .S1(n5921), .Q(
        n4990) );
  MUX41X1 U5955 ( .IN1(\FIFO[48][14] ), .IN3(\FIFO[50][14] ), .IN2(
        \FIFO[49][14] ), .IN4(\FIFO[51][14] ), .S0(n5827), .S1(n5921), .Q(
        n4991) );
  MUX41X1 U5956 ( .IN1(n4991), .IN3(n4989), .IN2(n4990), .IN4(n4988), .S0(
        n5744), .S1(n5763), .Q(n4992) );
  MUX41X1 U5957 ( .IN1(\FIFO[44][14] ), .IN3(\FIFO[46][14] ), .IN2(
        \FIFO[45][14] ), .IN4(\FIFO[47][14] ), .S0(n5827), .S1(n5921), .Q(
        n4993) );
  MUX41X1 U5958 ( .IN1(\FIFO[40][14] ), .IN3(\FIFO[42][14] ), .IN2(
        \FIFO[41][14] ), .IN4(\FIFO[43][14] ), .S0(n5827), .S1(n5921), .Q(
        n4994) );
  MUX41X1 U5959 ( .IN1(\FIFO[36][14] ), .IN3(\FIFO[38][14] ), .IN2(
        \FIFO[37][14] ), .IN4(\FIFO[39][14] ), .S0(n5827), .S1(n5921), .Q(
        n4995) );
  MUX41X1 U5960 ( .IN1(\FIFO[32][14] ), .IN3(\FIFO[34][14] ), .IN2(
        \FIFO[33][14] ), .IN4(\FIFO[35][14] ), .S0(n5827), .S1(n5921), .Q(
        n4996) );
  MUX41X1 U5961 ( .IN1(n4996), .IN3(n4994), .IN2(n4995), .IN4(n4993), .S0(
        n5744), .S1(n5763), .Q(n4997) );
  MUX41X1 U5962 ( .IN1(\FIFO[28][14] ), .IN3(\FIFO[30][14] ), .IN2(
        \FIFO[29][14] ), .IN4(\FIFO[31][14] ), .S0(n5828), .S1(n5922), .Q(
        n4998) );
  MUX41X1 U5963 ( .IN1(\FIFO[24][14] ), .IN3(\FIFO[26][14] ), .IN2(
        \FIFO[25][14] ), .IN4(\FIFO[27][14] ), .S0(n5828), .S1(n5922), .Q(
        n4999) );
  MUX41X1 U5964 ( .IN1(\FIFO[20][14] ), .IN3(\FIFO[22][14] ), .IN2(
        \FIFO[21][14] ), .IN4(\FIFO[23][14] ), .S0(n5828), .S1(n5922), .Q(
        n5000) );
  MUX41X1 U5965 ( .IN1(\FIFO[16][14] ), .IN3(\FIFO[18][14] ), .IN2(
        \FIFO[17][14] ), .IN4(\FIFO[19][14] ), .S0(n5828), .S1(n5922), .Q(
        n5001) );
  MUX41X1 U5966 ( .IN1(n5001), .IN3(n4999), .IN2(n5000), .IN4(n4998), .S0(
        n5744), .S1(n5763), .Q(n5002) );
  MUX41X1 U5967 ( .IN1(\FIFO[12][14] ), .IN3(\FIFO[14][14] ), .IN2(
        \FIFO[13][14] ), .IN4(\FIFO[15][14] ), .S0(n5828), .S1(n5922), .Q(
        n5003) );
  MUX41X1 U5968 ( .IN1(\FIFO[8][14] ), .IN3(\FIFO[10][14] ), .IN2(
        \FIFO[9][14] ), .IN4(\FIFO[11][14] ), .S0(n5828), .S1(n5922), .Q(n5004) );
  MUX41X1 U5969 ( .IN1(\FIFO[4][14] ), .IN3(\FIFO[6][14] ), .IN2(\FIFO[5][14] ), .IN4(\FIFO[7][14] ), .S0(n5828), .S1(n5922), .Q(n5005) );
  MUX41X1 U5970 ( .IN1(\FIFO[0][14] ), .IN3(\FIFO[2][14] ), .IN2(\FIFO[1][14] ), .IN4(\FIFO[3][14] ), .S0(n5828), .S1(n5922), .Q(n5006) );
  MUX41X1 U5971 ( .IN1(n5006), .IN3(n5004), .IN2(n5005), .IN4(n5003), .S0(
        n5744), .S1(n5763), .Q(n5007) );
  MUX41X1 U5972 ( .IN1(n5007), .IN3(n4997), .IN2(n5002), .IN4(n4992), .S0(
        n5728), .S1(n5732), .Q(n5008) );
  MUX21X1 U5973 ( .IN1(n5008), .IN2(n4987), .S(n5723), .Q(N236) );
  MUX41X1 U5974 ( .IN1(\FIFO[124][15] ), .IN3(\FIFO[126][15] ), .IN2(
        \FIFO[125][15] ), .IN4(\FIFO[127][15] ), .S0(n5828), .S1(n5922), .Q(
        n5009) );
  MUX41X1 U5975 ( .IN1(\FIFO[120][15] ), .IN3(\FIFO[122][15] ), .IN2(
        \FIFO[121][15] ), .IN4(\FIFO[123][15] ), .S0(n5828), .S1(n5922), .Q(
        n5010) );
  MUX41X1 U5976 ( .IN1(\FIFO[116][15] ), .IN3(\FIFO[118][15] ), .IN2(
        \FIFO[117][15] ), .IN4(\FIFO[119][15] ), .S0(n5828), .S1(n5922), .Q(
        n5011) );
  MUX41X1 U5977 ( .IN1(\FIFO[112][15] ), .IN3(\FIFO[114][15] ), .IN2(
        \FIFO[113][15] ), .IN4(\FIFO[115][15] ), .S0(n5828), .S1(n5922), .Q(
        n5012) );
  MUX41X1 U5978 ( .IN1(n5012), .IN3(n5010), .IN2(n5011), .IN4(n5009), .S0(
        n5744), .S1(n5763), .Q(n5013) );
  MUX41X1 U5979 ( .IN1(\FIFO[108][15] ), .IN3(\FIFO[110][15] ), .IN2(
        \FIFO[109][15] ), .IN4(\FIFO[111][15] ), .S0(n5829), .S1(n5923), .Q(
        n5014) );
  MUX41X1 U5980 ( .IN1(\FIFO[104][15] ), .IN3(\FIFO[106][15] ), .IN2(
        \FIFO[105][15] ), .IN4(\FIFO[107][15] ), .S0(n5829), .S1(n5923), .Q(
        n5015) );
  MUX41X1 U5981 ( .IN1(\FIFO[100][15] ), .IN3(\FIFO[102][15] ), .IN2(
        \FIFO[101][15] ), .IN4(\FIFO[103][15] ), .S0(n5829), .S1(n5923), .Q(
        n5016) );
  MUX41X1 U5982 ( .IN1(\FIFO[96][15] ), .IN3(\FIFO[98][15] ), .IN2(
        \FIFO[97][15] ), .IN4(\FIFO[99][15] ), .S0(n5829), .S1(n5923), .Q(
        n5017) );
  MUX41X1 U5983 ( .IN1(n5017), .IN3(n5015), .IN2(n5016), .IN4(n5014), .S0(
        n5744), .S1(n5763), .Q(n5018) );
  MUX41X1 U5984 ( .IN1(\FIFO[92][15] ), .IN3(\FIFO[94][15] ), .IN2(
        \FIFO[93][15] ), .IN4(\FIFO[95][15] ), .S0(n5829), .S1(n5923), .Q(
        n5019) );
  MUX41X1 U5985 ( .IN1(\FIFO[88][15] ), .IN3(\FIFO[90][15] ), .IN2(
        \FIFO[89][15] ), .IN4(\FIFO[91][15] ), .S0(n5829), .S1(n5923), .Q(
        n5020) );
  MUX41X1 U5986 ( .IN1(\FIFO[84][15] ), .IN3(\FIFO[86][15] ), .IN2(
        \FIFO[85][15] ), .IN4(\FIFO[87][15] ), .S0(n5829), .S1(n5923), .Q(
        n5021) );
  MUX41X1 U5987 ( .IN1(\FIFO[80][15] ), .IN3(\FIFO[82][15] ), .IN2(
        \FIFO[81][15] ), .IN4(\FIFO[83][15] ), .S0(n5829), .S1(n5923), .Q(
        n5022) );
  MUX41X1 U5988 ( .IN1(n5022), .IN3(n5020), .IN2(n5021), .IN4(n5019), .S0(
        n5744), .S1(n5763), .Q(n5023) );
  MUX41X1 U5989 ( .IN1(\FIFO[76][15] ), .IN3(\FIFO[78][15] ), .IN2(
        \FIFO[77][15] ), .IN4(\FIFO[79][15] ), .S0(n5829), .S1(n5923), .Q(
        n5024) );
  MUX41X1 U5990 ( .IN1(\FIFO[72][15] ), .IN3(\FIFO[74][15] ), .IN2(
        \FIFO[73][15] ), .IN4(\FIFO[75][15] ), .S0(n5829), .S1(n5923), .Q(
        n5025) );
  MUX41X1 U5991 ( .IN1(\FIFO[68][15] ), .IN3(\FIFO[70][15] ), .IN2(
        \FIFO[69][15] ), .IN4(\FIFO[71][15] ), .S0(n5829), .S1(n5923), .Q(
        n5026) );
  MUX41X1 U5992 ( .IN1(\FIFO[64][15] ), .IN3(\FIFO[66][15] ), .IN2(
        \FIFO[65][15] ), .IN4(\FIFO[67][15] ), .S0(n5829), .S1(n5923), .Q(
        n5027) );
  MUX41X1 U5993 ( .IN1(n5027), .IN3(n5025), .IN2(n5026), .IN4(n5024), .S0(
        n5744), .S1(n5763), .Q(n5028) );
  MUX41X1 U5994 ( .IN1(n5028), .IN3(n5018), .IN2(n5023), .IN4(n5013), .S0(
        n5728), .S1(n5732), .Q(n5029) );
  MUX41X1 U5995 ( .IN1(\FIFO[60][15] ), .IN3(\FIFO[62][15] ), .IN2(
        \FIFO[61][15] ), .IN4(\FIFO[63][15] ), .S0(n5830), .S1(n5924), .Q(
        n5030) );
  MUX41X1 U5996 ( .IN1(\FIFO[56][15] ), .IN3(\FIFO[58][15] ), .IN2(
        \FIFO[57][15] ), .IN4(\FIFO[59][15] ), .S0(n5830), .S1(n5924), .Q(
        n5031) );
  MUX41X1 U5997 ( .IN1(\FIFO[52][15] ), .IN3(\FIFO[54][15] ), .IN2(
        \FIFO[53][15] ), .IN4(\FIFO[55][15] ), .S0(n5830), .S1(n5924), .Q(
        n5032) );
  MUX41X1 U5998 ( .IN1(\FIFO[48][15] ), .IN3(\FIFO[50][15] ), .IN2(
        \FIFO[49][15] ), .IN4(\FIFO[51][15] ), .S0(n5830), .S1(n5924), .Q(
        n5033) );
  MUX41X1 U5999 ( .IN1(n5033), .IN3(n5031), .IN2(n5032), .IN4(n5030), .S0(
        n5745), .S1(n5764), .Q(n5034) );
  MUX41X1 U6000 ( .IN1(\FIFO[44][15] ), .IN3(\FIFO[46][15] ), .IN2(
        \FIFO[45][15] ), .IN4(\FIFO[47][15] ), .S0(n5830), .S1(n5924), .Q(
        n5035) );
  MUX41X1 U6001 ( .IN1(\FIFO[40][15] ), .IN3(\FIFO[42][15] ), .IN2(
        \FIFO[41][15] ), .IN4(\FIFO[43][15] ), .S0(n5830), .S1(n5924), .Q(
        n5036) );
  MUX41X1 U6002 ( .IN1(\FIFO[36][15] ), .IN3(\FIFO[38][15] ), .IN2(
        \FIFO[37][15] ), .IN4(\FIFO[39][15] ), .S0(n5830), .S1(n5924), .Q(
        n5037) );
  MUX41X1 U6003 ( .IN1(\FIFO[32][15] ), .IN3(\FIFO[34][15] ), .IN2(
        \FIFO[33][15] ), .IN4(\FIFO[35][15] ), .S0(n5830), .S1(n5924), .Q(
        n5038) );
  MUX41X1 U6004 ( .IN1(n5038), .IN3(n5036), .IN2(n5037), .IN4(n5035), .S0(
        n5745), .S1(n5764), .Q(n5039) );
  MUX41X1 U6005 ( .IN1(\FIFO[28][15] ), .IN3(\FIFO[30][15] ), .IN2(
        \FIFO[29][15] ), .IN4(\FIFO[31][15] ), .S0(n5830), .S1(n5924), .Q(
        n5040) );
  MUX41X1 U6006 ( .IN1(\FIFO[24][15] ), .IN3(\FIFO[26][15] ), .IN2(
        \FIFO[25][15] ), .IN4(\FIFO[27][15] ), .S0(n5830), .S1(n5924), .Q(
        n5041) );
  MUX41X1 U6007 ( .IN1(\FIFO[20][15] ), .IN3(\FIFO[22][15] ), .IN2(
        \FIFO[21][15] ), .IN4(\FIFO[23][15] ), .S0(n5830), .S1(n5924), .Q(
        n5042) );
  MUX41X1 U6008 ( .IN1(\FIFO[16][15] ), .IN3(\FIFO[18][15] ), .IN2(
        \FIFO[17][15] ), .IN4(\FIFO[19][15] ), .S0(n5830), .S1(n5924), .Q(
        n5043) );
  MUX41X1 U6009 ( .IN1(n5043), .IN3(n5041), .IN2(n5042), .IN4(n5040), .S0(
        n5745), .S1(n5764), .Q(n5044) );
  MUX41X1 U6010 ( .IN1(\FIFO[12][15] ), .IN3(\FIFO[14][15] ), .IN2(
        \FIFO[13][15] ), .IN4(\FIFO[15][15] ), .S0(n5831), .S1(n5925), .Q(
        n5045) );
  MUX41X1 U6011 ( .IN1(\FIFO[8][15] ), .IN3(\FIFO[10][15] ), .IN2(
        \FIFO[9][15] ), .IN4(\FIFO[11][15] ), .S0(n5831), .S1(n5925), .Q(n5046) );
  MUX41X1 U6012 ( .IN1(\FIFO[4][15] ), .IN3(\FIFO[6][15] ), .IN2(\FIFO[5][15] ), .IN4(\FIFO[7][15] ), .S0(n5831), .S1(n5925), .Q(n5047) );
  MUX41X1 U6013 ( .IN1(\FIFO[0][15] ), .IN3(\FIFO[2][15] ), .IN2(\FIFO[1][15] ), .IN4(\FIFO[3][15] ), .S0(n5831), .S1(n5925), .Q(n5048) );
  MUX41X1 U6014 ( .IN1(n5048), .IN3(n5046), .IN2(n5047), .IN4(n5045), .S0(
        n5745), .S1(n5764), .Q(n5049) );
  MUX41X1 U6015 ( .IN1(n5049), .IN3(n5039), .IN2(n5044), .IN4(n5034), .S0(
        n5728), .S1(n5732), .Q(n5050) );
  MUX21X1 U6016 ( .IN1(n5050), .IN2(n5029), .S(n5723), .Q(N235) );
  MUX41X1 U6017 ( .IN1(\FIFO[124][16] ), .IN3(\FIFO[126][16] ), .IN2(
        \FIFO[125][16] ), .IN4(\FIFO[127][16] ), .S0(n5831), .S1(n5925), .Q(
        n5051) );
  MUX41X1 U6018 ( .IN1(\FIFO[120][16] ), .IN3(\FIFO[122][16] ), .IN2(
        \FIFO[121][16] ), .IN4(\FIFO[123][16] ), .S0(n5831), .S1(n5925), .Q(
        n5052) );
  MUX41X1 U6019 ( .IN1(\FIFO[116][16] ), .IN3(\FIFO[118][16] ), .IN2(
        \FIFO[117][16] ), .IN4(\FIFO[119][16] ), .S0(n5831), .S1(n5925), .Q(
        n5053) );
  MUX41X1 U6020 ( .IN1(\FIFO[112][16] ), .IN3(\FIFO[114][16] ), .IN2(
        \FIFO[113][16] ), .IN4(\FIFO[115][16] ), .S0(n5831), .S1(n5925), .Q(
        n5054) );
  MUX41X1 U6021 ( .IN1(n5054), .IN3(n5052), .IN2(n5053), .IN4(n5051), .S0(
        n5745), .S1(n5764), .Q(n5055) );
  MUX41X1 U6022 ( .IN1(\FIFO[108][16] ), .IN3(\FIFO[110][16] ), .IN2(
        \FIFO[109][16] ), .IN4(\FIFO[111][16] ), .S0(n5831), .S1(n5925), .Q(
        n5056) );
  MUX41X1 U6023 ( .IN1(\FIFO[104][16] ), .IN3(\FIFO[106][16] ), .IN2(
        \FIFO[105][16] ), .IN4(\FIFO[107][16] ), .S0(n5831), .S1(n5925), .Q(
        n5057) );
  MUX41X1 U6024 ( .IN1(\FIFO[100][16] ), .IN3(\FIFO[102][16] ), .IN2(
        \FIFO[101][16] ), .IN4(\FIFO[103][16] ), .S0(n5831), .S1(n5925), .Q(
        n5058) );
  MUX41X1 U6025 ( .IN1(\FIFO[96][16] ), .IN3(\FIFO[98][16] ), .IN2(
        \FIFO[97][16] ), .IN4(\FIFO[99][16] ), .S0(n5831), .S1(n5925), .Q(
        n5059) );
  MUX41X1 U6026 ( .IN1(n5059), .IN3(n5057), .IN2(n5058), .IN4(n5056), .S0(
        n5745), .S1(n5764), .Q(n5060) );
  MUX41X1 U6027 ( .IN1(\FIFO[92][16] ), .IN3(\FIFO[94][16] ), .IN2(
        \FIFO[93][16] ), .IN4(\FIFO[95][16] ), .S0(n5832), .S1(n5926), .Q(
        n5061) );
  MUX41X1 U6028 ( .IN1(\FIFO[88][16] ), .IN3(\FIFO[90][16] ), .IN2(
        \FIFO[89][16] ), .IN4(\FIFO[91][16] ), .S0(n5832), .S1(n5926), .Q(
        n5062) );
  MUX41X1 U6029 ( .IN1(\FIFO[84][16] ), .IN3(\FIFO[86][16] ), .IN2(
        \FIFO[85][16] ), .IN4(\FIFO[87][16] ), .S0(n5832), .S1(n5926), .Q(
        n5063) );
  MUX41X1 U6030 ( .IN1(\FIFO[80][16] ), .IN3(\FIFO[82][16] ), .IN2(
        \FIFO[81][16] ), .IN4(\FIFO[83][16] ), .S0(n5832), .S1(n5926), .Q(
        n5064) );
  MUX41X1 U6031 ( .IN1(n5064), .IN3(n5062), .IN2(n5063), .IN4(n5061), .S0(
        n5745), .S1(n5764), .Q(n5065) );
  MUX41X1 U6032 ( .IN1(\FIFO[76][16] ), .IN3(\FIFO[78][16] ), .IN2(
        \FIFO[77][16] ), .IN4(\FIFO[79][16] ), .S0(n5832), .S1(n5926), .Q(
        n5066) );
  MUX41X1 U6033 ( .IN1(\FIFO[72][16] ), .IN3(\FIFO[74][16] ), .IN2(
        \FIFO[73][16] ), .IN4(\FIFO[75][16] ), .S0(n5832), .S1(n5926), .Q(
        n5067) );
  MUX41X1 U6034 ( .IN1(\FIFO[68][16] ), .IN3(\FIFO[70][16] ), .IN2(
        \FIFO[69][16] ), .IN4(\FIFO[71][16] ), .S0(n5832), .S1(n5926), .Q(
        n5068) );
  MUX41X1 U6035 ( .IN1(\FIFO[64][16] ), .IN3(\FIFO[66][16] ), .IN2(
        \FIFO[65][16] ), .IN4(\FIFO[67][16] ), .S0(n5832), .S1(n5926), .Q(
        n5069) );
  MUX41X1 U6036 ( .IN1(n5069), .IN3(n5067), .IN2(n5068), .IN4(n5066), .S0(
        n5745), .S1(n5764), .Q(n5070) );
  MUX41X1 U6037 ( .IN1(n5070), .IN3(n5060), .IN2(n5065), .IN4(n5055), .S0(
        n5728), .S1(n5732), .Q(n5071) );
  MUX41X1 U6038 ( .IN1(\FIFO[60][16] ), .IN3(\FIFO[62][16] ), .IN2(
        \FIFO[61][16] ), .IN4(\FIFO[63][16] ), .S0(n5832), .S1(n5926), .Q(
        n5072) );
  MUX41X1 U6039 ( .IN1(\FIFO[56][16] ), .IN3(\FIFO[58][16] ), .IN2(
        \FIFO[57][16] ), .IN4(\FIFO[59][16] ), .S0(n5832), .S1(n5926), .Q(
        n5073) );
  MUX41X1 U6040 ( .IN1(\FIFO[52][16] ), .IN3(\FIFO[54][16] ), .IN2(
        \FIFO[53][16] ), .IN4(\FIFO[55][16] ), .S0(n5832), .S1(n5926), .Q(
        n5074) );
  MUX41X1 U6041 ( .IN1(\FIFO[48][16] ), .IN3(\FIFO[50][16] ), .IN2(
        \FIFO[49][16] ), .IN4(\FIFO[51][16] ), .S0(n5832), .S1(n5926), .Q(
        n5075) );
  MUX41X1 U6042 ( .IN1(n5075), .IN3(n5073), .IN2(n5074), .IN4(n5072), .S0(
        n5745), .S1(n5764), .Q(n5076) );
  MUX41X1 U6043 ( .IN1(\FIFO[44][16] ), .IN3(\FIFO[46][16] ), .IN2(
        \FIFO[45][16] ), .IN4(\FIFO[47][16] ), .S0(n5833), .S1(n5927), .Q(
        n5077) );
  MUX41X1 U6044 ( .IN1(\FIFO[40][16] ), .IN3(\FIFO[42][16] ), .IN2(
        \FIFO[41][16] ), .IN4(\FIFO[43][16] ), .S0(n5833), .S1(n5927), .Q(
        n5078) );
  MUX41X1 U6045 ( .IN1(\FIFO[36][16] ), .IN3(\FIFO[38][16] ), .IN2(
        \FIFO[37][16] ), .IN4(\FIFO[39][16] ), .S0(n5833), .S1(n5927), .Q(
        n5079) );
  MUX41X1 U6046 ( .IN1(\FIFO[32][16] ), .IN3(\FIFO[34][16] ), .IN2(
        \FIFO[33][16] ), .IN4(\FIFO[35][16] ), .S0(n5833), .S1(n5927), .Q(
        n5080) );
  MUX41X1 U6047 ( .IN1(n5080), .IN3(n5078), .IN2(n5079), .IN4(n5077), .S0(
        n5745), .S1(n5764), .Q(n5081) );
  MUX41X1 U6048 ( .IN1(\FIFO[28][16] ), .IN3(\FIFO[30][16] ), .IN2(
        \FIFO[29][16] ), .IN4(\FIFO[31][16] ), .S0(n5833), .S1(n5927), .Q(
        n5082) );
  MUX41X1 U6049 ( .IN1(\FIFO[24][16] ), .IN3(\FIFO[26][16] ), .IN2(
        \FIFO[25][16] ), .IN4(\FIFO[27][16] ), .S0(n5833), .S1(n5927), .Q(
        n5083) );
  MUX41X1 U6050 ( .IN1(\FIFO[20][16] ), .IN3(\FIFO[22][16] ), .IN2(
        \FIFO[21][16] ), .IN4(\FIFO[23][16] ), .S0(n5833), .S1(n5927), .Q(
        n5084) );
  MUX41X1 U6051 ( .IN1(\FIFO[16][16] ), .IN3(\FIFO[18][16] ), .IN2(
        \FIFO[17][16] ), .IN4(\FIFO[19][16] ), .S0(n5833), .S1(n5927), .Q(
        n5085) );
  MUX41X1 U6052 ( .IN1(n5085), .IN3(n5083), .IN2(n5084), .IN4(n5082), .S0(
        n5745), .S1(n5764), .Q(n5086) );
  MUX41X1 U6053 ( .IN1(\FIFO[12][16] ), .IN3(\FIFO[14][16] ), .IN2(
        \FIFO[13][16] ), .IN4(\FIFO[15][16] ), .S0(n5833), .S1(n5927), .Q(
        n5087) );
  MUX41X1 U6054 ( .IN1(\FIFO[8][16] ), .IN3(\FIFO[10][16] ), .IN2(
        \FIFO[9][16] ), .IN4(\FIFO[11][16] ), .S0(n5833), .S1(n5927), .Q(n5088) );
  MUX41X1 U6055 ( .IN1(\FIFO[4][16] ), .IN3(\FIFO[6][16] ), .IN2(\FIFO[5][16] ), .IN4(\FIFO[7][16] ), .S0(n5833), .S1(n5927), .Q(n5089) );
  MUX41X1 U6056 ( .IN1(\FIFO[0][16] ), .IN3(\FIFO[2][16] ), .IN2(\FIFO[1][16] ), .IN4(\FIFO[3][16] ), .S0(n5833), .S1(n5927), .Q(n5090) );
  MUX41X1 U6057 ( .IN1(n5090), .IN3(n5088), .IN2(n5089), .IN4(n5087), .S0(
        n5745), .S1(n5764), .Q(n5091) );
  MUX41X1 U6058 ( .IN1(n5091), .IN3(n5081), .IN2(n5086), .IN4(n5076), .S0(
        n5728), .S1(n5732), .Q(n5092) );
  MUX21X1 U6059 ( .IN1(n5092), .IN2(n5071), .S(n5723), .Q(N234) );
  MUX41X1 U6060 ( .IN1(\FIFO[124][17] ), .IN3(\FIFO[126][17] ), .IN2(
        \FIFO[125][17] ), .IN4(\FIFO[127][17] ), .S0(n5834), .S1(n5928), .Q(
        n5093) );
  MUX41X1 U6061 ( .IN1(\FIFO[120][17] ), .IN3(\FIFO[122][17] ), .IN2(
        \FIFO[121][17] ), .IN4(\FIFO[123][17] ), .S0(n5834), .S1(n5928), .Q(
        n5094) );
  MUX41X1 U6062 ( .IN1(\FIFO[116][17] ), .IN3(\FIFO[118][17] ), .IN2(
        \FIFO[117][17] ), .IN4(\FIFO[119][17] ), .S0(n5834), .S1(n5928), .Q(
        n5095) );
  MUX41X1 U6063 ( .IN1(\FIFO[112][17] ), .IN3(\FIFO[114][17] ), .IN2(
        \FIFO[113][17] ), .IN4(\FIFO[115][17] ), .S0(n5834), .S1(n5928), .Q(
        n5096) );
  MUX41X1 U6064 ( .IN1(n5096), .IN3(n5094), .IN2(n5095), .IN4(n5093), .S0(
        n5746), .S1(n5765), .Q(n5097) );
  MUX41X1 U6065 ( .IN1(\FIFO[108][17] ), .IN3(\FIFO[110][17] ), .IN2(
        \FIFO[109][17] ), .IN4(\FIFO[111][17] ), .S0(n5834), .S1(n5928), .Q(
        n5098) );
  MUX41X1 U6066 ( .IN1(\FIFO[104][17] ), .IN3(\FIFO[106][17] ), .IN2(
        \FIFO[105][17] ), .IN4(\FIFO[107][17] ), .S0(n5834), .S1(n5928), .Q(
        n5099) );
  MUX41X1 U6067 ( .IN1(\FIFO[100][17] ), .IN3(\FIFO[102][17] ), .IN2(
        \FIFO[101][17] ), .IN4(\FIFO[103][17] ), .S0(n5834), .S1(n5928), .Q(
        n5100) );
  MUX41X1 U6068 ( .IN1(\FIFO[96][17] ), .IN3(\FIFO[98][17] ), .IN2(
        \FIFO[97][17] ), .IN4(\FIFO[99][17] ), .S0(n5834), .S1(n5928), .Q(
        n5101) );
  MUX41X1 U6069 ( .IN1(n5101), .IN3(n5099), .IN2(n5100), .IN4(n5098), .S0(
        n5746), .S1(n5765), .Q(n5102) );
  MUX41X1 U6070 ( .IN1(\FIFO[92][17] ), .IN3(\FIFO[94][17] ), .IN2(
        \FIFO[93][17] ), .IN4(\FIFO[95][17] ), .S0(n5834), .S1(n5928), .Q(
        n5103) );
  MUX41X1 U6071 ( .IN1(\FIFO[88][17] ), .IN3(\FIFO[90][17] ), .IN2(
        \FIFO[89][17] ), .IN4(\FIFO[91][17] ), .S0(n5834), .S1(n5928), .Q(
        n5104) );
  MUX41X1 U6072 ( .IN1(\FIFO[84][17] ), .IN3(\FIFO[86][17] ), .IN2(
        \FIFO[85][17] ), .IN4(\FIFO[87][17] ), .S0(n5834), .S1(n5928), .Q(
        n5105) );
  MUX41X1 U6073 ( .IN1(\FIFO[80][17] ), .IN3(\FIFO[82][17] ), .IN2(
        \FIFO[81][17] ), .IN4(\FIFO[83][17] ), .S0(n5834), .S1(n5928), .Q(
        n5106) );
  MUX41X1 U6074 ( .IN1(n5106), .IN3(n5104), .IN2(n5105), .IN4(n5103), .S0(
        n5746), .S1(n5765), .Q(n5107) );
  MUX41X1 U6075 ( .IN1(\FIFO[76][17] ), .IN3(\FIFO[78][17] ), .IN2(
        \FIFO[77][17] ), .IN4(\FIFO[79][17] ), .S0(n5835), .S1(n5929), .Q(
        n5108) );
  MUX41X1 U6076 ( .IN1(\FIFO[72][17] ), .IN3(\FIFO[74][17] ), .IN2(
        \FIFO[73][17] ), .IN4(\FIFO[75][17] ), .S0(n5835), .S1(n5929), .Q(
        n5109) );
  MUX41X1 U6077 ( .IN1(\FIFO[68][17] ), .IN3(\FIFO[70][17] ), .IN2(
        \FIFO[69][17] ), .IN4(\FIFO[71][17] ), .S0(n5835), .S1(n5929), .Q(
        n5110) );
  MUX41X1 U6078 ( .IN1(\FIFO[64][17] ), .IN3(\FIFO[66][17] ), .IN2(
        \FIFO[65][17] ), .IN4(\FIFO[67][17] ), .S0(n5835), .S1(n5929), .Q(
        n5111) );
  MUX41X1 U6079 ( .IN1(n5111), .IN3(n5109), .IN2(n5110), .IN4(n5108), .S0(
        n5746), .S1(n5765), .Q(n5112) );
  MUX41X1 U6080 ( .IN1(n5112), .IN3(n5102), .IN2(n5107), .IN4(n5097), .S0(
        n5728), .S1(n5732), .Q(n5113) );
  MUX41X1 U6081 ( .IN1(\FIFO[60][17] ), .IN3(\FIFO[62][17] ), .IN2(
        \FIFO[61][17] ), .IN4(\FIFO[63][17] ), .S0(n5835), .S1(n5929), .Q(
        n5114) );
  MUX41X1 U6082 ( .IN1(\FIFO[56][17] ), .IN3(\FIFO[58][17] ), .IN2(
        \FIFO[57][17] ), .IN4(\FIFO[59][17] ), .S0(n5835), .S1(n5929), .Q(
        n5115) );
  MUX41X1 U6083 ( .IN1(\FIFO[52][17] ), .IN3(\FIFO[54][17] ), .IN2(
        \FIFO[53][17] ), .IN4(\FIFO[55][17] ), .S0(n5835), .S1(n5929), .Q(
        n5116) );
  MUX41X1 U6084 ( .IN1(\FIFO[48][17] ), .IN3(\FIFO[50][17] ), .IN2(
        \FIFO[49][17] ), .IN4(\FIFO[51][17] ), .S0(n5835), .S1(n5929), .Q(
        n5117) );
  MUX41X1 U6085 ( .IN1(n5117), .IN3(n5115), .IN2(n5116), .IN4(n5114), .S0(
        n5746), .S1(n5765), .Q(n5118) );
  MUX41X1 U6086 ( .IN1(\FIFO[44][17] ), .IN3(\FIFO[46][17] ), .IN2(
        \FIFO[45][17] ), .IN4(\FIFO[47][17] ), .S0(n5835), .S1(n5929), .Q(
        n5119) );
  MUX41X1 U6087 ( .IN1(\FIFO[40][17] ), .IN3(\FIFO[42][17] ), .IN2(
        \FIFO[41][17] ), .IN4(\FIFO[43][17] ), .S0(n5835), .S1(n5929), .Q(
        n5120) );
  MUX41X1 U6088 ( .IN1(\FIFO[36][17] ), .IN3(\FIFO[38][17] ), .IN2(
        \FIFO[37][17] ), .IN4(\FIFO[39][17] ), .S0(n5835), .S1(n5929), .Q(
        n5121) );
  MUX41X1 U6089 ( .IN1(\FIFO[32][17] ), .IN3(\FIFO[34][17] ), .IN2(
        \FIFO[33][17] ), .IN4(\FIFO[35][17] ), .S0(n5835), .S1(n5929), .Q(
        n5122) );
  MUX41X1 U6090 ( .IN1(n5122), .IN3(n5120), .IN2(n5121), .IN4(n5119), .S0(
        n5746), .S1(n5765), .Q(n5123) );
  MUX41X1 U6091 ( .IN1(\FIFO[28][17] ), .IN3(\FIFO[30][17] ), .IN2(
        \FIFO[29][17] ), .IN4(\FIFO[31][17] ), .S0(n5836), .S1(n5930), .Q(
        n5124) );
  MUX41X1 U6092 ( .IN1(\FIFO[24][17] ), .IN3(\FIFO[26][17] ), .IN2(
        \FIFO[25][17] ), .IN4(\FIFO[27][17] ), .S0(n5836), .S1(n5930), .Q(
        n5125) );
  MUX41X1 U6093 ( .IN1(\FIFO[20][17] ), .IN3(\FIFO[22][17] ), .IN2(
        \FIFO[21][17] ), .IN4(\FIFO[23][17] ), .S0(n5836), .S1(n5930), .Q(
        n5126) );
  MUX41X1 U6094 ( .IN1(\FIFO[16][17] ), .IN3(\FIFO[18][17] ), .IN2(
        \FIFO[17][17] ), .IN4(\FIFO[19][17] ), .S0(n5836), .S1(n5930), .Q(
        n5127) );
  MUX41X1 U6095 ( .IN1(n5127), .IN3(n5125), .IN2(n5126), .IN4(n5124), .S0(
        n5746), .S1(n5765), .Q(n5128) );
  MUX41X1 U6096 ( .IN1(\FIFO[12][17] ), .IN3(\FIFO[14][17] ), .IN2(
        \FIFO[13][17] ), .IN4(\FIFO[15][17] ), .S0(n5836), .S1(n5930), .Q(
        n5129) );
  MUX41X1 U6097 ( .IN1(\FIFO[8][17] ), .IN3(\FIFO[10][17] ), .IN2(
        \FIFO[9][17] ), .IN4(\FIFO[11][17] ), .S0(n5836), .S1(n5930), .Q(n5130) );
  MUX41X1 U6098 ( .IN1(\FIFO[4][17] ), .IN3(\FIFO[6][17] ), .IN2(\FIFO[5][17] ), .IN4(\FIFO[7][17] ), .S0(n5836), .S1(n5930), .Q(n5131) );
  MUX41X1 U6099 ( .IN1(\FIFO[0][17] ), .IN3(\FIFO[2][17] ), .IN2(\FIFO[1][17] ), .IN4(\FIFO[3][17] ), .S0(n5836), .S1(n5930), .Q(n5132) );
  MUX41X1 U6100 ( .IN1(n5132), .IN3(n5130), .IN2(n5131), .IN4(n5129), .S0(
        n5746), .S1(n5765), .Q(n5133) );
  MUX41X1 U6101 ( .IN1(n5133), .IN3(n5123), .IN2(n5128), .IN4(n5118), .S0(
        n5728), .S1(n5732), .Q(n5134) );
  MUX21X1 U6102 ( .IN1(n5134), .IN2(n5113), .S(n5723), .Q(N233) );
  MUX41X1 U6103 ( .IN1(\FIFO[124][18] ), .IN3(\FIFO[126][18] ), .IN2(
        \FIFO[125][18] ), .IN4(\FIFO[127][18] ), .S0(n5836), .S1(n5930), .Q(
        n5135) );
  MUX41X1 U6104 ( .IN1(\FIFO[120][18] ), .IN3(\FIFO[122][18] ), .IN2(
        \FIFO[121][18] ), .IN4(\FIFO[123][18] ), .S0(n5836), .S1(n5930), .Q(
        n5136) );
  MUX41X1 U6105 ( .IN1(\FIFO[116][18] ), .IN3(\FIFO[118][18] ), .IN2(
        \FIFO[117][18] ), .IN4(\FIFO[119][18] ), .S0(n5836), .S1(n5930), .Q(
        n5137) );
  MUX41X1 U6106 ( .IN1(\FIFO[112][18] ), .IN3(\FIFO[114][18] ), .IN2(
        \FIFO[113][18] ), .IN4(\FIFO[115][18] ), .S0(n5836), .S1(n5930), .Q(
        n5138) );
  MUX41X1 U6107 ( .IN1(n5138), .IN3(n5136), .IN2(n5137), .IN4(n5135), .S0(
        n5746), .S1(n5765), .Q(n5139) );
  MUX41X1 U6108 ( .IN1(\FIFO[108][18] ), .IN3(\FIFO[110][18] ), .IN2(
        \FIFO[109][18] ), .IN4(\FIFO[111][18] ), .S0(n5837), .S1(n5931), .Q(
        n5140) );
  MUX41X1 U6109 ( .IN1(\FIFO[104][18] ), .IN3(\FIFO[106][18] ), .IN2(
        \FIFO[105][18] ), .IN4(\FIFO[107][18] ), .S0(n5837), .S1(n5931), .Q(
        n5141) );
  MUX41X1 U6110 ( .IN1(\FIFO[100][18] ), .IN3(\FIFO[102][18] ), .IN2(
        \FIFO[101][18] ), .IN4(\FIFO[103][18] ), .S0(n5837), .S1(n5931), .Q(
        n5142) );
  MUX41X1 U6111 ( .IN1(\FIFO[96][18] ), .IN3(\FIFO[98][18] ), .IN2(
        \FIFO[97][18] ), .IN4(\FIFO[99][18] ), .S0(n5837), .S1(n5931), .Q(
        n5143) );
  MUX41X1 U6112 ( .IN1(n5143), .IN3(n5141), .IN2(n5142), .IN4(n5140), .S0(
        n5746), .S1(n5765), .Q(n5144) );
  MUX41X1 U6113 ( .IN1(\FIFO[92][18] ), .IN3(\FIFO[94][18] ), .IN2(
        \FIFO[93][18] ), .IN4(\FIFO[95][18] ), .S0(n5837), .S1(n5931), .Q(
        n5145) );
  MUX41X1 U6114 ( .IN1(\FIFO[88][18] ), .IN3(\FIFO[90][18] ), .IN2(
        \FIFO[89][18] ), .IN4(\FIFO[91][18] ), .S0(n5837), .S1(n5931), .Q(
        n5146) );
  MUX41X1 U6115 ( .IN1(\FIFO[84][18] ), .IN3(\FIFO[86][18] ), .IN2(
        \FIFO[85][18] ), .IN4(\FIFO[87][18] ), .S0(n5837), .S1(n5931), .Q(
        n5147) );
  MUX41X1 U6116 ( .IN1(\FIFO[80][18] ), .IN3(\FIFO[82][18] ), .IN2(
        \FIFO[81][18] ), .IN4(\FIFO[83][18] ), .S0(n5837), .S1(n5931), .Q(
        n5148) );
  MUX41X1 U6117 ( .IN1(n5148), .IN3(n5146), .IN2(n5147), .IN4(n5145), .S0(
        n5746), .S1(n5765), .Q(n5149) );
  MUX41X1 U6118 ( .IN1(\FIFO[76][18] ), .IN3(\FIFO[78][18] ), .IN2(
        \FIFO[77][18] ), .IN4(\FIFO[79][18] ), .S0(n5837), .S1(n5931), .Q(
        n5150) );
  MUX41X1 U6119 ( .IN1(\FIFO[72][18] ), .IN3(\FIFO[74][18] ), .IN2(
        \FIFO[73][18] ), .IN4(\FIFO[75][18] ), .S0(n5837), .S1(n5931), .Q(
        n5151) );
  MUX41X1 U6120 ( .IN1(\FIFO[68][18] ), .IN3(\FIFO[70][18] ), .IN2(
        \FIFO[69][18] ), .IN4(\FIFO[71][18] ), .S0(n5837), .S1(n5931), .Q(
        n5152) );
  MUX41X1 U6121 ( .IN1(\FIFO[64][18] ), .IN3(\FIFO[66][18] ), .IN2(
        \FIFO[65][18] ), .IN4(\FIFO[67][18] ), .S0(n5837), .S1(n5931), .Q(
        n5153) );
  MUX41X1 U6122 ( .IN1(n5153), .IN3(n5151), .IN2(n5152), .IN4(n5150), .S0(
        n5746), .S1(n5765), .Q(n5154) );
  MUX41X1 U6123 ( .IN1(n5154), .IN3(n5144), .IN2(n5149), .IN4(n5139), .S0(
        n5728), .S1(n5732), .Q(n5155) );
  MUX41X1 U6124 ( .IN1(\FIFO[60][18] ), .IN3(\FIFO[62][18] ), .IN2(
        \FIFO[61][18] ), .IN4(\FIFO[63][18] ), .S0(n5838), .S1(n5932), .Q(
        n5156) );
  MUX41X1 U6125 ( .IN1(\FIFO[56][18] ), .IN3(\FIFO[58][18] ), .IN2(
        \FIFO[57][18] ), .IN4(\FIFO[59][18] ), .S0(n5838), .S1(n5932), .Q(
        n5157) );
  MUX41X1 U6126 ( .IN1(\FIFO[52][18] ), .IN3(\FIFO[54][18] ), .IN2(
        \FIFO[53][18] ), .IN4(\FIFO[55][18] ), .S0(n5838), .S1(n5932), .Q(
        n5158) );
  MUX41X1 U6127 ( .IN1(\FIFO[48][18] ), .IN3(\FIFO[50][18] ), .IN2(
        \FIFO[49][18] ), .IN4(\FIFO[51][18] ), .S0(n5838), .S1(n5932), .Q(
        n5159) );
  MUX41X1 U6128 ( .IN1(n5159), .IN3(n5157), .IN2(n5158), .IN4(n5156), .S0(
        n5747), .S1(n5766), .Q(n5160) );
  MUX41X1 U6129 ( .IN1(\FIFO[44][18] ), .IN3(\FIFO[46][18] ), .IN2(
        \FIFO[45][18] ), .IN4(\FIFO[47][18] ), .S0(n5838), .S1(n5932), .Q(
        n5161) );
  MUX41X1 U6130 ( .IN1(\FIFO[40][18] ), .IN3(\FIFO[42][18] ), .IN2(
        \FIFO[41][18] ), .IN4(\FIFO[43][18] ), .S0(n5838), .S1(n5932), .Q(
        n5162) );
  MUX41X1 U6131 ( .IN1(\FIFO[36][18] ), .IN3(\FIFO[38][18] ), .IN2(
        \FIFO[37][18] ), .IN4(\FIFO[39][18] ), .S0(n5838), .S1(n5932), .Q(
        n5163) );
  MUX41X1 U6132 ( .IN1(\FIFO[32][18] ), .IN3(\FIFO[34][18] ), .IN2(
        \FIFO[33][18] ), .IN4(\FIFO[35][18] ), .S0(n5838), .S1(n5932), .Q(
        n5164) );
  MUX41X1 U6133 ( .IN1(n5164), .IN3(n5162), .IN2(n5163), .IN4(n5161), .S0(
        n5747), .S1(n5766), .Q(n5165) );
  MUX41X1 U6134 ( .IN1(\FIFO[28][18] ), .IN3(\FIFO[30][18] ), .IN2(
        \FIFO[29][18] ), .IN4(\FIFO[31][18] ), .S0(n5838), .S1(n5932), .Q(
        n5166) );
  MUX41X1 U6135 ( .IN1(\FIFO[24][18] ), .IN3(\FIFO[26][18] ), .IN2(
        \FIFO[25][18] ), .IN4(\FIFO[27][18] ), .S0(n5838), .S1(n5932), .Q(
        n5167) );
  MUX41X1 U6136 ( .IN1(\FIFO[20][18] ), .IN3(\FIFO[22][18] ), .IN2(
        \FIFO[21][18] ), .IN4(\FIFO[23][18] ), .S0(n5838), .S1(n5932), .Q(
        n5168) );
  MUX41X1 U6137 ( .IN1(\FIFO[16][18] ), .IN3(\FIFO[18][18] ), .IN2(
        \FIFO[17][18] ), .IN4(\FIFO[19][18] ), .S0(n5838), .S1(n5932), .Q(
        n5169) );
  MUX41X1 U6138 ( .IN1(n5169), .IN3(n5167), .IN2(n5168), .IN4(n5166), .S0(
        n5747), .S1(n5766), .Q(n5170) );
  MUX41X1 U6139 ( .IN1(\FIFO[12][18] ), .IN3(\FIFO[14][18] ), .IN2(
        \FIFO[13][18] ), .IN4(\FIFO[15][18] ), .S0(n5839), .S1(n5933), .Q(
        n5171) );
  MUX41X1 U6140 ( .IN1(\FIFO[8][18] ), .IN3(\FIFO[10][18] ), .IN2(
        \FIFO[9][18] ), .IN4(\FIFO[11][18] ), .S0(n5839), .S1(n5933), .Q(n5172) );
  MUX41X1 U6141 ( .IN1(\FIFO[4][18] ), .IN3(\FIFO[6][18] ), .IN2(\FIFO[5][18] ), .IN4(\FIFO[7][18] ), .S0(n5839), .S1(n5933), .Q(n5173) );
  MUX41X1 U6142 ( .IN1(\FIFO[0][18] ), .IN3(\FIFO[2][18] ), .IN2(\FIFO[1][18] ), .IN4(\FIFO[3][18] ), .S0(n5839), .S1(n5933), .Q(n5174) );
  MUX41X1 U6143 ( .IN1(n5174), .IN3(n5172), .IN2(n5173), .IN4(n5171), .S0(
        n5747), .S1(n5766), .Q(n5175) );
  MUX41X1 U6144 ( .IN1(n5175), .IN3(n5165), .IN2(n5170), .IN4(n5160), .S0(
        n5728), .S1(n5732), .Q(n5176) );
  MUX21X1 U6145 ( .IN1(n5176), .IN2(n5155), .S(n5723), .Q(N232) );
  MUX41X1 U6146 ( .IN1(\FIFO[124][19] ), .IN3(\FIFO[126][19] ), .IN2(
        \FIFO[125][19] ), .IN4(\FIFO[127][19] ), .S0(n5839), .S1(n5933), .Q(
        n5177) );
  MUX41X1 U6147 ( .IN1(\FIFO[120][19] ), .IN3(\FIFO[122][19] ), .IN2(
        \FIFO[121][19] ), .IN4(\FIFO[123][19] ), .S0(n5839), .S1(n5933), .Q(
        n5178) );
  MUX41X1 U6148 ( .IN1(\FIFO[116][19] ), .IN3(\FIFO[118][19] ), .IN2(
        \FIFO[117][19] ), .IN4(\FIFO[119][19] ), .S0(n5839), .S1(n5933), .Q(
        n5179) );
  MUX41X1 U6149 ( .IN1(\FIFO[112][19] ), .IN3(\FIFO[114][19] ), .IN2(
        \FIFO[113][19] ), .IN4(\FIFO[115][19] ), .S0(n5839), .S1(n5933), .Q(
        n5180) );
  MUX41X1 U6150 ( .IN1(n5180), .IN3(n5178), .IN2(n5179), .IN4(n5177), .S0(
        n5747), .S1(n5766), .Q(n5181) );
  MUX41X1 U6151 ( .IN1(\FIFO[108][19] ), .IN3(\FIFO[110][19] ), .IN2(
        \FIFO[109][19] ), .IN4(\FIFO[111][19] ), .S0(n5839), .S1(n5933), .Q(
        n5182) );
  MUX41X1 U6152 ( .IN1(\FIFO[104][19] ), .IN3(\FIFO[106][19] ), .IN2(
        \FIFO[105][19] ), .IN4(\FIFO[107][19] ), .S0(n5839), .S1(n5933), .Q(
        n5183) );
  MUX41X1 U6153 ( .IN1(\FIFO[100][19] ), .IN3(\FIFO[102][19] ), .IN2(
        \FIFO[101][19] ), .IN4(\FIFO[103][19] ), .S0(n5839), .S1(n5933), .Q(
        n5184) );
  MUX41X1 U6154 ( .IN1(\FIFO[96][19] ), .IN3(\FIFO[98][19] ), .IN2(
        \FIFO[97][19] ), .IN4(\FIFO[99][19] ), .S0(n5839), .S1(n5933), .Q(
        n5185) );
  MUX41X1 U6155 ( .IN1(n5185), .IN3(n5183), .IN2(n5184), .IN4(n5182), .S0(
        n5747), .S1(n5766), .Q(n5186) );
  MUX41X1 U6156 ( .IN1(\FIFO[92][19] ), .IN3(\FIFO[94][19] ), .IN2(
        \FIFO[93][19] ), .IN4(\FIFO[95][19] ), .S0(n5840), .S1(n5934), .Q(
        n5187) );
  MUX41X1 U6157 ( .IN1(\FIFO[88][19] ), .IN3(\FIFO[90][19] ), .IN2(
        \FIFO[89][19] ), .IN4(\FIFO[91][19] ), .S0(n5840), .S1(n5934), .Q(
        n5188) );
  MUX41X1 U6158 ( .IN1(\FIFO[84][19] ), .IN3(\FIFO[86][19] ), .IN2(
        \FIFO[85][19] ), .IN4(\FIFO[87][19] ), .S0(n5840), .S1(n5934), .Q(
        n5189) );
  MUX41X1 U6159 ( .IN1(\FIFO[80][19] ), .IN3(\FIFO[82][19] ), .IN2(
        \FIFO[81][19] ), .IN4(\FIFO[83][19] ), .S0(n5840), .S1(n5934), .Q(
        n5190) );
  MUX41X1 U6160 ( .IN1(n5190), .IN3(n5188), .IN2(n5189), .IN4(n5187), .S0(
        n5747), .S1(n5766), .Q(n5191) );
  MUX41X1 U6161 ( .IN1(\FIFO[76][19] ), .IN3(\FIFO[78][19] ), .IN2(
        \FIFO[77][19] ), .IN4(\FIFO[79][19] ), .S0(n5840), .S1(n5934), .Q(
        n5192) );
  MUX41X1 U6162 ( .IN1(\FIFO[72][19] ), .IN3(\FIFO[74][19] ), .IN2(
        \FIFO[73][19] ), .IN4(\FIFO[75][19] ), .S0(n5840), .S1(n5934), .Q(
        n5193) );
  MUX41X1 U6163 ( .IN1(\FIFO[68][19] ), .IN3(\FIFO[70][19] ), .IN2(
        \FIFO[69][19] ), .IN4(\FIFO[71][19] ), .S0(n5840), .S1(n5934), .Q(
        n5194) );
  MUX41X1 U6164 ( .IN1(\FIFO[64][19] ), .IN3(\FIFO[66][19] ), .IN2(
        \FIFO[65][19] ), .IN4(\FIFO[67][19] ), .S0(n5840), .S1(n5934), .Q(
        n5195) );
  MUX41X1 U6165 ( .IN1(n5195), .IN3(n5193), .IN2(n5194), .IN4(n5192), .S0(
        n5747), .S1(n5766), .Q(n5196) );
  MUX41X1 U6166 ( .IN1(n5196), .IN3(n5186), .IN2(n5191), .IN4(n5181), .S0(
        n5728), .S1(n5732), .Q(n5197) );
  MUX41X1 U6167 ( .IN1(\FIFO[60][19] ), .IN3(\FIFO[62][19] ), .IN2(
        \FIFO[61][19] ), .IN4(\FIFO[63][19] ), .S0(n5840), .S1(n5934), .Q(
        n5198) );
  MUX41X1 U6168 ( .IN1(\FIFO[56][19] ), .IN3(\FIFO[58][19] ), .IN2(
        \FIFO[57][19] ), .IN4(\FIFO[59][19] ), .S0(n5840), .S1(n5934), .Q(
        n5199) );
  MUX41X1 U6169 ( .IN1(\FIFO[52][19] ), .IN3(\FIFO[54][19] ), .IN2(
        \FIFO[53][19] ), .IN4(\FIFO[55][19] ), .S0(n5840), .S1(n5934), .Q(
        n5200) );
  MUX41X1 U6170 ( .IN1(\FIFO[48][19] ), .IN3(\FIFO[50][19] ), .IN2(
        \FIFO[49][19] ), .IN4(\FIFO[51][19] ), .S0(n5840), .S1(n5934), .Q(
        n5201) );
  MUX41X1 U6171 ( .IN1(n5201), .IN3(n5199), .IN2(n5200), .IN4(n5198), .S0(
        n5747), .S1(n5766), .Q(n5202) );
  MUX41X1 U6172 ( .IN1(\FIFO[44][19] ), .IN3(\FIFO[46][19] ), .IN2(
        \FIFO[45][19] ), .IN4(\FIFO[47][19] ), .S0(n5841), .S1(n5935), .Q(
        n5203) );
  MUX41X1 U6173 ( .IN1(\FIFO[40][19] ), .IN3(\FIFO[42][19] ), .IN2(
        \FIFO[41][19] ), .IN4(\FIFO[43][19] ), .S0(n5841), .S1(n5935), .Q(
        n5204) );
  MUX41X1 U6174 ( .IN1(\FIFO[36][19] ), .IN3(\FIFO[38][19] ), .IN2(
        \FIFO[37][19] ), .IN4(\FIFO[39][19] ), .S0(n5841), .S1(n5935), .Q(
        n5205) );
  MUX41X1 U6175 ( .IN1(\FIFO[32][19] ), .IN3(\FIFO[34][19] ), .IN2(
        \FIFO[33][19] ), .IN4(\FIFO[35][19] ), .S0(n5841), .S1(n5935), .Q(
        n5206) );
  MUX41X1 U6176 ( .IN1(n5206), .IN3(n5204), .IN2(n5205), .IN4(n5203), .S0(
        n5747), .S1(n5766), .Q(n5207) );
  MUX41X1 U6177 ( .IN1(\FIFO[28][19] ), .IN3(\FIFO[30][19] ), .IN2(
        \FIFO[29][19] ), .IN4(\FIFO[31][19] ), .S0(n5841), .S1(n5935), .Q(
        n5208) );
  MUX41X1 U6178 ( .IN1(\FIFO[24][19] ), .IN3(\FIFO[26][19] ), .IN2(
        \FIFO[25][19] ), .IN4(\FIFO[27][19] ), .S0(n5841), .S1(n5935), .Q(
        n5209) );
  MUX41X1 U6179 ( .IN1(\FIFO[20][19] ), .IN3(\FIFO[22][19] ), .IN2(
        \FIFO[21][19] ), .IN4(\FIFO[23][19] ), .S0(n5841), .S1(n5935), .Q(
        n5210) );
  MUX41X1 U6180 ( .IN1(\FIFO[16][19] ), .IN3(\FIFO[18][19] ), .IN2(
        \FIFO[17][19] ), .IN4(\FIFO[19][19] ), .S0(n5841), .S1(n5935), .Q(
        n5211) );
  MUX41X1 U6181 ( .IN1(n5211), .IN3(n5209), .IN2(n5210), .IN4(n5208), .S0(
        n5747), .S1(n5766), .Q(n5212) );
  MUX41X1 U6182 ( .IN1(\FIFO[12][19] ), .IN3(\FIFO[14][19] ), .IN2(
        \FIFO[13][19] ), .IN4(\FIFO[15][19] ), .S0(n5841), .S1(n5935), .Q(
        n5213) );
  MUX41X1 U6183 ( .IN1(\FIFO[8][19] ), .IN3(\FIFO[10][19] ), .IN2(
        \FIFO[9][19] ), .IN4(\FIFO[11][19] ), .S0(n5841), .S1(n5935), .Q(n5214) );
  MUX41X1 U6184 ( .IN1(\FIFO[4][19] ), .IN3(\FIFO[6][19] ), .IN2(\FIFO[5][19] ), .IN4(\FIFO[7][19] ), .S0(n5841), .S1(n5935), .Q(n5215) );
  MUX41X1 U6185 ( .IN1(\FIFO[0][19] ), .IN3(\FIFO[2][19] ), .IN2(\FIFO[1][19] ), .IN4(\FIFO[3][19] ), .S0(n5841), .S1(n5935), .Q(n5216) );
  MUX41X1 U6186 ( .IN1(n5216), .IN3(n5214), .IN2(n5215), .IN4(n5213), .S0(
        n5747), .S1(n5766), .Q(n5217) );
  MUX41X1 U6187 ( .IN1(n5217), .IN3(n5207), .IN2(n5212), .IN4(n5202), .S0(
        n5728), .S1(n5732), .Q(n5218) );
  MUX21X1 U6188 ( .IN1(n5218), .IN2(n5197), .S(n5723), .Q(N231) );
  MUX41X1 U6189 ( .IN1(\FIFO[124][20] ), .IN3(\FIFO[126][20] ), .IN2(
        \FIFO[125][20] ), .IN4(\FIFO[127][20] ), .S0(n5842), .S1(n5936), .Q(
        n5219) );
  MUX41X1 U6190 ( .IN1(\FIFO[120][20] ), .IN3(\FIFO[122][20] ), .IN2(
        \FIFO[121][20] ), .IN4(\FIFO[123][20] ), .S0(n5842), .S1(n5936), .Q(
        n5220) );
  MUX41X1 U6191 ( .IN1(\FIFO[116][20] ), .IN3(\FIFO[118][20] ), .IN2(
        \FIFO[117][20] ), .IN4(\FIFO[119][20] ), .S0(n5842), .S1(n5936), .Q(
        n5221) );
  MUX41X1 U6192 ( .IN1(\FIFO[112][20] ), .IN3(\FIFO[114][20] ), .IN2(
        \FIFO[113][20] ), .IN4(\FIFO[115][20] ), .S0(n5842), .S1(n5936), .Q(
        n5222) );
  MUX41X1 U6193 ( .IN1(n5222), .IN3(n5220), .IN2(n5221), .IN4(n5219), .S0(
        n5748), .S1(n5767), .Q(n5223) );
  MUX41X1 U6194 ( .IN1(\FIFO[108][20] ), .IN3(\FIFO[110][20] ), .IN2(
        \FIFO[109][20] ), .IN4(\FIFO[111][20] ), .S0(n5842), .S1(n5936), .Q(
        n5224) );
  MUX41X1 U6195 ( .IN1(\FIFO[104][20] ), .IN3(\FIFO[106][20] ), .IN2(
        \FIFO[105][20] ), .IN4(\FIFO[107][20] ), .S0(n5842), .S1(n5936), .Q(
        n5225) );
  MUX41X1 U6196 ( .IN1(\FIFO[100][20] ), .IN3(\FIFO[102][20] ), .IN2(
        \FIFO[101][20] ), .IN4(\FIFO[103][20] ), .S0(n5842), .S1(n5936), .Q(
        n5226) );
  MUX41X1 U6197 ( .IN1(\FIFO[96][20] ), .IN3(\FIFO[98][20] ), .IN2(
        \FIFO[97][20] ), .IN4(\FIFO[99][20] ), .S0(n5842), .S1(n5936), .Q(
        n5227) );
  MUX41X1 U6198 ( .IN1(n5227), .IN3(n5225), .IN2(n5226), .IN4(n5224), .S0(
        n5748), .S1(n5767), .Q(n5228) );
  MUX41X1 U6199 ( .IN1(\FIFO[92][20] ), .IN3(\FIFO[94][20] ), .IN2(
        \FIFO[93][20] ), .IN4(\FIFO[95][20] ), .S0(n5842), .S1(n5936), .Q(
        n5229) );
  MUX41X1 U6200 ( .IN1(\FIFO[88][20] ), .IN3(\FIFO[90][20] ), .IN2(
        \FIFO[89][20] ), .IN4(\FIFO[91][20] ), .S0(n5842), .S1(n5936), .Q(
        n5230) );
  MUX41X1 U6201 ( .IN1(\FIFO[84][20] ), .IN3(\FIFO[86][20] ), .IN2(
        \FIFO[85][20] ), .IN4(\FIFO[87][20] ), .S0(n5842), .S1(n5936), .Q(
        n5231) );
  MUX41X1 U6202 ( .IN1(\FIFO[80][20] ), .IN3(\FIFO[82][20] ), .IN2(
        \FIFO[81][20] ), .IN4(\FIFO[83][20] ), .S0(n5842), .S1(n5936), .Q(
        n5232) );
  MUX41X1 U6203 ( .IN1(n5232), .IN3(n5230), .IN2(n5231), .IN4(n5229), .S0(
        n5748), .S1(n5767), .Q(n5233) );
  MUX41X1 U6204 ( .IN1(\FIFO[76][20] ), .IN3(\FIFO[78][20] ), .IN2(
        \FIFO[77][20] ), .IN4(\FIFO[79][20] ), .S0(n5843), .S1(n5937), .Q(
        n5234) );
  MUX41X1 U6205 ( .IN1(\FIFO[72][20] ), .IN3(\FIFO[74][20] ), .IN2(
        \FIFO[73][20] ), .IN4(\FIFO[75][20] ), .S0(n5843), .S1(n5937), .Q(
        n5235) );
  MUX41X1 U6206 ( .IN1(\FIFO[68][20] ), .IN3(\FIFO[70][20] ), .IN2(
        \FIFO[69][20] ), .IN4(\FIFO[71][20] ), .S0(n5843), .S1(n5937), .Q(
        n5236) );
  MUX41X1 U6207 ( .IN1(\FIFO[64][20] ), .IN3(\FIFO[66][20] ), .IN2(
        \FIFO[65][20] ), .IN4(\FIFO[67][20] ), .S0(n5843), .S1(n5937), .Q(
        n5237) );
  MUX41X1 U6208 ( .IN1(n5237), .IN3(n5235), .IN2(n5236), .IN4(n5234), .S0(
        n5748), .S1(n5767), .Q(n5238) );
  MUX41X1 U6209 ( .IN1(n5238), .IN3(n5228), .IN2(n5233), .IN4(n5223), .S0(
        n5729), .S1(n5733), .Q(n5239) );
  MUX41X1 U6210 ( .IN1(\FIFO[60][20] ), .IN3(\FIFO[62][20] ), .IN2(
        \FIFO[61][20] ), .IN4(\FIFO[63][20] ), .S0(n5843), .S1(n5937), .Q(
        n5240) );
  MUX41X1 U6211 ( .IN1(\FIFO[56][20] ), .IN3(\FIFO[58][20] ), .IN2(
        \FIFO[57][20] ), .IN4(\FIFO[59][20] ), .S0(n5843), .S1(n5937), .Q(
        n5241) );
  MUX41X1 U6212 ( .IN1(\FIFO[52][20] ), .IN3(\FIFO[54][20] ), .IN2(
        \FIFO[53][20] ), .IN4(\FIFO[55][20] ), .S0(n5843), .S1(n5937), .Q(
        n5242) );
  MUX41X1 U6213 ( .IN1(\FIFO[48][20] ), .IN3(\FIFO[50][20] ), .IN2(
        \FIFO[49][20] ), .IN4(\FIFO[51][20] ), .S0(n5843), .S1(n5937), .Q(
        n5243) );
  MUX41X1 U6214 ( .IN1(n5243), .IN3(n5241), .IN2(n5242), .IN4(n5240), .S0(
        n5748), .S1(n5767), .Q(n5244) );
  MUX41X1 U6215 ( .IN1(\FIFO[44][20] ), .IN3(\FIFO[46][20] ), .IN2(
        \FIFO[45][20] ), .IN4(\FIFO[47][20] ), .S0(n5843), .S1(n5937), .Q(
        n5245) );
  MUX41X1 U6216 ( .IN1(\FIFO[40][20] ), .IN3(\FIFO[42][20] ), .IN2(
        \FIFO[41][20] ), .IN4(\FIFO[43][20] ), .S0(n5843), .S1(n5937), .Q(
        n5246) );
  MUX41X1 U6217 ( .IN1(\FIFO[36][20] ), .IN3(\FIFO[38][20] ), .IN2(
        \FIFO[37][20] ), .IN4(\FIFO[39][20] ), .S0(n5843), .S1(n5937), .Q(
        n5247) );
  MUX41X1 U6218 ( .IN1(\FIFO[32][20] ), .IN3(\FIFO[34][20] ), .IN2(
        \FIFO[33][20] ), .IN4(\FIFO[35][20] ), .S0(n5843), .S1(n5937), .Q(
        n5248) );
  MUX41X1 U6219 ( .IN1(n5248), .IN3(n5246), .IN2(n5247), .IN4(n5245), .S0(
        n5748), .S1(n5767), .Q(n5249) );
  MUX41X1 U6220 ( .IN1(\FIFO[28][20] ), .IN3(\FIFO[30][20] ), .IN2(
        \FIFO[29][20] ), .IN4(\FIFO[31][20] ), .S0(n5844), .S1(n5938), .Q(
        n5250) );
  MUX41X1 U6221 ( .IN1(\FIFO[24][20] ), .IN3(\FIFO[26][20] ), .IN2(
        \FIFO[25][20] ), .IN4(\FIFO[27][20] ), .S0(n5844), .S1(n5938), .Q(
        n5251) );
  MUX41X1 U6222 ( .IN1(\FIFO[20][20] ), .IN3(\FIFO[22][20] ), .IN2(
        \FIFO[21][20] ), .IN4(\FIFO[23][20] ), .S0(n5844), .S1(n5938), .Q(
        n5252) );
  MUX41X1 U6223 ( .IN1(\FIFO[16][20] ), .IN3(\FIFO[18][20] ), .IN2(
        \FIFO[17][20] ), .IN4(\FIFO[19][20] ), .S0(n5844), .S1(n5938), .Q(
        n5253) );
  MUX41X1 U6224 ( .IN1(n5253), .IN3(n5251), .IN2(n5252), .IN4(n5250), .S0(
        n5748), .S1(n5767), .Q(n5254) );
  MUX41X1 U6225 ( .IN1(\FIFO[12][20] ), .IN3(\FIFO[14][20] ), .IN2(
        \FIFO[13][20] ), .IN4(\FIFO[15][20] ), .S0(n5844), .S1(n5938), .Q(
        n5255) );
  MUX41X1 U6226 ( .IN1(\FIFO[8][20] ), .IN3(\FIFO[10][20] ), .IN2(
        \FIFO[9][20] ), .IN4(\FIFO[11][20] ), .S0(n5844), .S1(n5938), .Q(n5256) );
  MUX41X1 U6227 ( .IN1(\FIFO[4][20] ), .IN3(\FIFO[6][20] ), .IN2(\FIFO[5][20] ), .IN4(\FIFO[7][20] ), .S0(n5844), .S1(n5938), .Q(n5257) );
  MUX41X1 U6228 ( .IN1(\FIFO[0][20] ), .IN3(\FIFO[2][20] ), .IN2(\FIFO[1][20] ), .IN4(\FIFO[3][20] ), .S0(n5844), .S1(n5938), .Q(n5258) );
  MUX41X1 U6229 ( .IN1(n5258), .IN3(n5256), .IN2(n5257), .IN4(n5255), .S0(
        n5748), .S1(n5767), .Q(n5259) );
  MUX41X1 U6230 ( .IN1(n5259), .IN3(n5249), .IN2(n5254), .IN4(n5244), .S0(
        n5729), .S1(n5733), .Q(n5260) );
  MUX21X1 U6231 ( .IN1(n5260), .IN2(n5239), .S(n5724), .Q(N230) );
  MUX41X1 U6232 ( .IN1(\FIFO[124][21] ), .IN3(\FIFO[126][21] ), .IN2(
        \FIFO[125][21] ), .IN4(\FIFO[127][21] ), .S0(n5844), .S1(n5938), .Q(
        n5261) );
  MUX41X1 U6233 ( .IN1(\FIFO[120][21] ), .IN3(\FIFO[122][21] ), .IN2(
        \FIFO[121][21] ), .IN4(\FIFO[123][21] ), .S0(n5844), .S1(n5938), .Q(
        n5262) );
  MUX41X1 U6234 ( .IN1(\FIFO[116][21] ), .IN3(\FIFO[118][21] ), .IN2(
        \FIFO[117][21] ), .IN4(\FIFO[119][21] ), .S0(n5844), .S1(n5938), .Q(
        n5263) );
  MUX41X1 U6235 ( .IN1(\FIFO[112][21] ), .IN3(\FIFO[114][21] ), .IN2(
        \FIFO[113][21] ), .IN4(\FIFO[115][21] ), .S0(n5844), .S1(n5938), .Q(
        n5264) );
  MUX41X1 U6236 ( .IN1(n5264), .IN3(n5262), .IN2(n5263), .IN4(n5261), .S0(
        n5748), .S1(n5767), .Q(n5265) );
  MUX41X1 U6237 ( .IN1(\FIFO[108][21] ), .IN3(\FIFO[110][21] ), .IN2(
        \FIFO[109][21] ), .IN4(\FIFO[111][21] ), .S0(n5845), .S1(n5939), .Q(
        n5266) );
  MUX41X1 U6238 ( .IN1(\FIFO[104][21] ), .IN3(\FIFO[106][21] ), .IN2(
        \FIFO[105][21] ), .IN4(\FIFO[107][21] ), .S0(n5845), .S1(n5939), .Q(
        n5267) );
  MUX41X1 U6239 ( .IN1(\FIFO[100][21] ), .IN3(\FIFO[102][21] ), .IN2(
        \FIFO[101][21] ), .IN4(\FIFO[103][21] ), .S0(n5845), .S1(n5939), .Q(
        n5268) );
  MUX41X1 U6240 ( .IN1(\FIFO[96][21] ), .IN3(\FIFO[98][21] ), .IN2(
        \FIFO[97][21] ), .IN4(\FIFO[99][21] ), .S0(n5845), .S1(n5939), .Q(
        n5269) );
  MUX41X1 U6241 ( .IN1(n5269), .IN3(n5267), .IN2(n5268), .IN4(n5266), .S0(
        n5748), .S1(n5767), .Q(n5270) );
  MUX41X1 U6242 ( .IN1(\FIFO[92][21] ), .IN3(\FIFO[94][21] ), .IN2(
        \FIFO[93][21] ), .IN4(\FIFO[95][21] ), .S0(n5845), .S1(n5939), .Q(
        n5271) );
  MUX41X1 U6243 ( .IN1(\FIFO[88][21] ), .IN3(\FIFO[90][21] ), .IN2(
        \FIFO[89][21] ), .IN4(\FIFO[91][21] ), .S0(n5845), .S1(n5939), .Q(
        n5272) );
  MUX41X1 U6244 ( .IN1(\FIFO[84][21] ), .IN3(\FIFO[86][21] ), .IN2(
        \FIFO[85][21] ), .IN4(\FIFO[87][21] ), .S0(n5845), .S1(n5939), .Q(
        n5273) );
  MUX41X1 U6245 ( .IN1(\FIFO[80][21] ), .IN3(\FIFO[82][21] ), .IN2(
        \FIFO[81][21] ), .IN4(\FIFO[83][21] ), .S0(n5845), .S1(n5939), .Q(
        n5274) );
  MUX41X1 U6246 ( .IN1(n5274), .IN3(n5272), .IN2(n5273), .IN4(n5271), .S0(
        n5748), .S1(n5767), .Q(n5275) );
  MUX41X1 U6247 ( .IN1(\FIFO[76][21] ), .IN3(\FIFO[78][21] ), .IN2(
        \FIFO[77][21] ), .IN4(\FIFO[79][21] ), .S0(n5845), .S1(n5939), .Q(
        n5276) );
  MUX41X1 U6248 ( .IN1(\FIFO[72][21] ), .IN3(\FIFO[74][21] ), .IN2(
        \FIFO[73][21] ), .IN4(\FIFO[75][21] ), .S0(n5845), .S1(n5939), .Q(
        n5277) );
  MUX41X1 U6249 ( .IN1(\FIFO[68][21] ), .IN3(\FIFO[70][21] ), .IN2(
        \FIFO[69][21] ), .IN4(\FIFO[71][21] ), .S0(n5845), .S1(n5939), .Q(
        n5278) );
  MUX41X1 U6250 ( .IN1(\FIFO[64][21] ), .IN3(\FIFO[66][21] ), .IN2(
        \FIFO[65][21] ), .IN4(\FIFO[67][21] ), .S0(n5845), .S1(n5939), .Q(
        n5279) );
  MUX41X1 U6251 ( .IN1(n5279), .IN3(n5277), .IN2(n5278), .IN4(n5276), .S0(
        n5748), .S1(n5767), .Q(n5280) );
  MUX41X1 U6252 ( .IN1(n5280), .IN3(n5270), .IN2(n5275), .IN4(n5265), .S0(
        n5729), .S1(n5733), .Q(n5281) );
  MUX41X1 U6253 ( .IN1(\FIFO[60][21] ), .IN3(\FIFO[62][21] ), .IN2(
        \FIFO[61][21] ), .IN4(\FIFO[63][21] ), .S0(n5846), .S1(n5940), .Q(
        n5282) );
  MUX41X1 U6254 ( .IN1(\FIFO[56][21] ), .IN3(\FIFO[58][21] ), .IN2(
        \FIFO[57][21] ), .IN4(\FIFO[59][21] ), .S0(n5846), .S1(n5940), .Q(
        n5283) );
  MUX41X1 U6255 ( .IN1(\FIFO[52][21] ), .IN3(\FIFO[54][21] ), .IN2(
        \FIFO[53][21] ), .IN4(\FIFO[55][21] ), .S0(n5846), .S1(n5940), .Q(
        n5284) );
  MUX41X1 U6256 ( .IN1(\FIFO[48][21] ), .IN3(\FIFO[50][21] ), .IN2(
        \FIFO[49][21] ), .IN4(\FIFO[51][21] ), .S0(n5846), .S1(n5940), .Q(
        n5285) );
  MUX41X1 U6257 ( .IN1(n5285), .IN3(n5283), .IN2(n5284), .IN4(n5282), .S0(
        n5749), .S1(n5768), .Q(n5286) );
  MUX41X1 U6258 ( .IN1(\FIFO[44][21] ), .IN3(\FIFO[46][21] ), .IN2(
        \FIFO[45][21] ), .IN4(\FIFO[47][21] ), .S0(n5846), .S1(n5940), .Q(
        n5287) );
  MUX41X1 U6259 ( .IN1(\FIFO[40][21] ), .IN3(\FIFO[42][21] ), .IN2(
        \FIFO[41][21] ), .IN4(\FIFO[43][21] ), .S0(n5846), .S1(n5940), .Q(
        n5288) );
  MUX41X1 U6260 ( .IN1(\FIFO[36][21] ), .IN3(\FIFO[38][21] ), .IN2(
        \FIFO[37][21] ), .IN4(\FIFO[39][21] ), .S0(n5846), .S1(n5940), .Q(
        n5289) );
  MUX41X1 U6261 ( .IN1(\FIFO[32][21] ), .IN3(\FIFO[34][21] ), .IN2(
        \FIFO[33][21] ), .IN4(\FIFO[35][21] ), .S0(n5846), .S1(n5940), .Q(
        n5290) );
  MUX41X1 U6262 ( .IN1(n5290), .IN3(n5288), .IN2(n5289), .IN4(n5287), .S0(
        n5749), .S1(n5768), .Q(n5291) );
  MUX41X1 U6263 ( .IN1(\FIFO[28][21] ), .IN3(\FIFO[30][21] ), .IN2(
        \FIFO[29][21] ), .IN4(\FIFO[31][21] ), .S0(n5846), .S1(n5940), .Q(
        n5292) );
  MUX41X1 U6264 ( .IN1(\FIFO[24][21] ), .IN3(\FIFO[26][21] ), .IN2(
        \FIFO[25][21] ), .IN4(\FIFO[27][21] ), .S0(n5846), .S1(n5940), .Q(
        n5293) );
  MUX41X1 U6265 ( .IN1(\FIFO[20][21] ), .IN3(\FIFO[22][21] ), .IN2(
        \FIFO[21][21] ), .IN4(\FIFO[23][21] ), .S0(n5846), .S1(n5940), .Q(
        n5294) );
  MUX41X1 U6266 ( .IN1(\FIFO[16][21] ), .IN3(\FIFO[18][21] ), .IN2(
        \FIFO[17][21] ), .IN4(\FIFO[19][21] ), .S0(n5846), .S1(n5940), .Q(
        n5295) );
  MUX41X1 U6267 ( .IN1(n5295), .IN3(n5293), .IN2(n5294), .IN4(n5292), .S0(
        n5749), .S1(n5768), .Q(n5296) );
  MUX41X1 U6268 ( .IN1(\FIFO[12][21] ), .IN3(\FIFO[14][21] ), .IN2(
        \FIFO[13][21] ), .IN4(\FIFO[15][21] ), .S0(n5847), .S1(n5941), .Q(
        n5297) );
  MUX41X1 U6269 ( .IN1(\FIFO[8][21] ), .IN3(\FIFO[10][21] ), .IN2(
        \FIFO[9][21] ), .IN4(\FIFO[11][21] ), .S0(n5847), .S1(n5941), .Q(n5298) );
  MUX41X1 U6270 ( .IN1(\FIFO[4][21] ), .IN3(\FIFO[6][21] ), .IN2(\FIFO[5][21] ), .IN4(\FIFO[7][21] ), .S0(n5847), .S1(n5941), .Q(n5299) );
  MUX41X1 U6271 ( .IN1(\FIFO[0][21] ), .IN3(\FIFO[2][21] ), .IN2(\FIFO[1][21] ), .IN4(\FIFO[3][21] ), .S0(n5847), .S1(n5941), .Q(n5300) );
  MUX41X1 U6272 ( .IN1(n5300), .IN3(n5298), .IN2(n5299), .IN4(n5297), .S0(
        n5749), .S1(n5768), .Q(n5301) );
  MUX41X1 U6273 ( .IN1(n5301), .IN3(n5291), .IN2(n5296), .IN4(n5286), .S0(
        n5729), .S1(n5733), .Q(n5302) );
  MUX21X1 U6274 ( .IN1(n5302), .IN2(n5281), .S(n5724), .Q(N229) );
  MUX41X1 U6275 ( .IN1(\FIFO[124][22] ), .IN3(\FIFO[126][22] ), .IN2(
        \FIFO[125][22] ), .IN4(\FIFO[127][22] ), .S0(n5847), .S1(n5941), .Q(
        n5303) );
  MUX41X1 U6276 ( .IN1(\FIFO[120][22] ), .IN3(\FIFO[122][22] ), .IN2(
        \FIFO[121][22] ), .IN4(\FIFO[123][22] ), .S0(n5847), .S1(n5941), .Q(
        n5304) );
  MUX41X1 U6277 ( .IN1(\FIFO[116][22] ), .IN3(\FIFO[118][22] ), .IN2(
        \FIFO[117][22] ), .IN4(\FIFO[119][22] ), .S0(n5847), .S1(n5941), .Q(
        n5305) );
  MUX41X1 U6278 ( .IN1(\FIFO[112][22] ), .IN3(\FIFO[114][22] ), .IN2(
        \FIFO[113][22] ), .IN4(\FIFO[115][22] ), .S0(n5847), .S1(n5941), .Q(
        n5306) );
  MUX41X1 U6279 ( .IN1(n5306), .IN3(n5304), .IN2(n5305), .IN4(n5303), .S0(
        n5749), .S1(n5768), .Q(n5307) );
  MUX41X1 U6280 ( .IN1(\FIFO[108][22] ), .IN3(\FIFO[110][22] ), .IN2(
        \FIFO[109][22] ), .IN4(\FIFO[111][22] ), .S0(n5847), .S1(n5941), .Q(
        n5308) );
  MUX41X1 U6281 ( .IN1(\FIFO[104][22] ), .IN3(\FIFO[106][22] ), .IN2(
        \FIFO[105][22] ), .IN4(\FIFO[107][22] ), .S0(n5847), .S1(n5941), .Q(
        n5309) );
  MUX41X1 U6282 ( .IN1(\FIFO[100][22] ), .IN3(\FIFO[102][22] ), .IN2(
        \FIFO[101][22] ), .IN4(\FIFO[103][22] ), .S0(n5847), .S1(n5941), .Q(
        n5310) );
  MUX41X1 U6283 ( .IN1(\FIFO[96][22] ), .IN3(\FIFO[98][22] ), .IN2(
        \FIFO[97][22] ), .IN4(\FIFO[99][22] ), .S0(n5847), .S1(n5941), .Q(
        n5311) );
  MUX41X1 U6284 ( .IN1(n5311), .IN3(n5309), .IN2(n5310), .IN4(n5308), .S0(
        n5749), .S1(n5768), .Q(n5312) );
  MUX41X1 U6285 ( .IN1(\FIFO[92][22] ), .IN3(\FIFO[94][22] ), .IN2(
        \FIFO[93][22] ), .IN4(\FIFO[95][22] ), .S0(n5848), .S1(n5942), .Q(
        n5313) );
  MUX41X1 U6286 ( .IN1(\FIFO[88][22] ), .IN3(\FIFO[90][22] ), .IN2(
        \FIFO[89][22] ), .IN4(\FIFO[91][22] ), .S0(n5848), .S1(n5942), .Q(
        n5314) );
  MUX41X1 U6287 ( .IN1(\FIFO[84][22] ), .IN3(\FIFO[86][22] ), .IN2(
        \FIFO[85][22] ), .IN4(\FIFO[87][22] ), .S0(n5848), .S1(n5942), .Q(
        n5315) );
  MUX41X1 U6288 ( .IN1(\FIFO[80][22] ), .IN3(\FIFO[82][22] ), .IN2(
        \FIFO[81][22] ), .IN4(\FIFO[83][22] ), .S0(n5848), .S1(n5942), .Q(
        n5316) );
  MUX41X1 U6289 ( .IN1(n5316), .IN3(n5314), .IN2(n5315), .IN4(n5313), .S0(
        n5749), .S1(n5768), .Q(n5317) );
  MUX41X1 U6290 ( .IN1(\FIFO[76][22] ), .IN3(\FIFO[78][22] ), .IN2(
        \FIFO[77][22] ), .IN4(\FIFO[79][22] ), .S0(n5848), .S1(n5942), .Q(
        n5318) );
  MUX41X1 U6291 ( .IN1(\FIFO[72][22] ), .IN3(\FIFO[74][22] ), .IN2(
        \FIFO[73][22] ), .IN4(\FIFO[75][22] ), .S0(n5848), .S1(n5942), .Q(
        n5319) );
  MUX41X1 U6292 ( .IN1(\FIFO[68][22] ), .IN3(\FIFO[70][22] ), .IN2(
        \FIFO[69][22] ), .IN4(\FIFO[71][22] ), .S0(n5848), .S1(n5942), .Q(
        n5320) );
  MUX41X1 U6293 ( .IN1(\FIFO[64][22] ), .IN3(\FIFO[66][22] ), .IN2(
        \FIFO[65][22] ), .IN4(\FIFO[67][22] ), .S0(n5848), .S1(n5942), .Q(
        n5321) );
  MUX41X1 U6294 ( .IN1(n5321), .IN3(n5319), .IN2(n5320), .IN4(n5318), .S0(
        n5749), .S1(n5768), .Q(n5322) );
  MUX41X1 U6295 ( .IN1(n5322), .IN3(n5312), .IN2(n5317), .IN4(n5307), .S0(
        n5729), .S1(n5733), .Q(n5323) );
  MUX41X1 U6296 ( .IN1(\FIFO[60][22] ), .IN3(\FIFO[62][22] ), .IN2(
        \FIFO[61][22] ), .IN4(\FIFO[63][22] ), .S0(n5848), .S1(n5942), .Q(
        n5324) );
  MUX41X1 U6297 ( .IN1(\FIFO[56][22] ), .IN3(\FIFO[58][22] ), .IN2(
        \FIFO[57][22] ), .IN4(\FIFO[59][22] ), .S0(n5848), .S1(n5942), .Q(
        n5325) );
  MUX41X1 U6298 ( .IN1(\FIFO[52][22] ), .IN3(\FIFO[54][22] ), .IN2(
        \FIFO[53][22] ), .IN4(\FIFO[55][22] ), .S0(n5848), .S1(n5942), .Q(
        n5326) );
  MUX41X1 U6299 ( .IN1(\FIFO[48][22] ), .IN3(\FIFO[50][22] ), .IN2(
        \FIFO[49][22] ), .IN4(\FIFO[51][22] ), .S0(n5848), .S1(n5942), .Q(
        n5327) );
  MUX41X1 U6300 ( .IN1(n5327), .IN3(n5325), .IN2(n5326), .IN4(n5324), .S0(
        n5749), .S1(n5768), .Q(n5328) );
  MUX41X1 U6301 ( .IN1(\FIFO[44][22] ), .IN3(\FIFO[46][22] ), .IN2(
        \FIFO[45][22] ), .IN4(\FIFO[47][22] ), .S0(n5849), .S1(n5943), .Q(
        n5329) );
  MUX41X1 U6302 ( .IN1(\FIFO[40][22] ), .IN3(\FIFO[42][22] ), .IN2(
        \FIFO[41][22] ), .IN4(\FIFO[43][22] ), .S0(n5849), .S1(n5943), .Q(
        n5330) );
  MUX41X1 U6303 ( .IN1(\FIFO[36][22] ), .IN3(\FIFO[38][22] ), .IN2(
        \FIFO[37][22] ), .IN4(\FIFO[39][22] ), .S0(n5849), .S1(n5943), .Q(
        n5331) );
  MUX41X1 U6304 ( .IN1(\FIFO[32][22] ), .IN3(\FIFO[34][22] ), .IN2(
        \FIFO[33][22] ), .IN4(\FIFO[35][22] ), .S0(n5849), .S1(n5943), .Q(
        n5332) );
  MUX41X1 U6305 ( .IN1(n5332), .IN3(n5330), .IN2(n5331), .IN4(n5329), .S0(
        n5749), .S1(n5768), .Q(n5333) );
  MUX41X1 U6306 ( .IN1(\FIFO[28][22] ), .IN3(\FIFO[30][22] ), .IN2(
        \FIFO[29][22] ), .IN4(\FIFO[31][22] ), .S0(n5849), .S1(n5943), .Q(
        n5334) );
  MUX41X1 U6307 ( .IN1(\FIFO[24][22] ), .IN3(\FIFO[26][22] ), .IN2(
        \FIFO[25][22] ), .IN4(\FIFO[27][22] ), .S0(n5849), .S1(n5943), .Q(
        n5335) );
  MUX41X1 U6308 ( .IN1(\FIFO[20][22] ), .IN3(\FIFO[22][22] ), .IN2(
        \FIFO[21][22] ), .IN4(\FIFO[23][22] ), .S0(n5849), .S1(n5943), .Q(
        n5336) );
  MUX41X1 U6309 ( .IN1(\FIFO[16][22] ), .IN3(\FIFO[18][22] ), .IN2(
        \FIFO[17][22] ), .IN4(\FIFO[19][22] ), .S0(n5849), .S1(n5943), .Q(
        n5337) );
  MUX41X1 U6310 ( .IN1(n5337), .IN3(n5335), .IN2(n5336), .IN4(n5334), .S0(
        n5749), .S1(n5768), .Q(n5338) );
  MUX41X1 U6311 ( .IN1(\FIFO[12][22] ), .IN3(\FIFO[14][22] ), .IN2(
        \FIFO[13][22] ), .IN4(\FIFO[15][22] ), .S0(n5849), .S1(n5943), .Q(
        n5339) );
  MUX41X1 U6312 ( .IN1(\FIFO[8][22] ), .IN3(\FIFO[10][22] ), .IN2(
        \FIFO[9][22] ), .IN4(\FIFO[11][22] ), .S0(n5849), .S1(n5943), .Q(n5340) );
  MUX41X1 U6313 ( .IN1(\FIFO[4][22] ), .IN3(\FIFO[6][22] ), .IN2(\FIFO[5][22] ), .IN4(\FIFO[7][22] ), .S0(n5849), .S1(n5943), .Q(n5341) );
  MUX41X1 U6314 ( .IN1(\FIFO[0][22] ), .IN3(\FIFO[2][22] ), .IN2(\FIFO[1][22] ), .IN4(\FIFO[3][22] ), .S0(n5849), .S1(n5943), .Q(n5342) );
  MUX41X1 U6315 ( .IN1(n5342), .IN3(n5340), .IN2(n5341), .IN4(n5339), .S0(
        n5749), .S1(n5768), .Q(n5343) );
  MUX41X1 U6316 ( .IN1(n5343), .IN3(n5333), .IN2(n5338), .IN4(n5328), .S0(
        n5729), .S1(n5733), .Q(n5344) );
  MUX21X1 U6317 ( .IN1(n5344), .IN2(n5323), .S(n5724), .Q(N228) );
  MUX41X1 U6318 ( .IN1(\FIFO[124][23] ), .IN3(\FIFO[126][23] ), .IN2(
        \FIFO[125][23] ), .IN4(\FIFO[127][23] ), .S0(n5850), .S1(n5944), .Q(
        n5345) );
  MUX41X1 U6319 ( .IN1(\FIFO[120][23] ), .IN3(\FIFO[122][23] ), .IN2(
        \FIFO[121][23] ), .IN4(\FIFO[123][23] ), .S0(n5850), .S1(n5944), .Q(
        n5346) );
  MUX41X1 U6320 ( .IN1(\FIFO[116][23] ), .IN3(\FIFO[118][23] ), .IN2(
        \FIFO[117][23] ), .IN4(\FIFO[119][23] ), .S0(n5850), .S1(n5944), .Q(
        n5347) );
  MUX41X1 U6321 ( .IN1(\FIFO[112][23] ), .IN3(\FIFO[114][23] ), .IN2(
        \FIFO[113][23] ), .IN4(\FIFO[115][23] ), .S0(n5850), .S1(n5944), .Q(
        n5348) );
  MUX41X1 U6322 ( .IN1(n5348), .IN3(n5346), .IN2(n5347), .IN4(n5345), .S0(
        n5750), .S1(n5769), .Q(n5349) );
  MUX41X1 U6323 ( .IN1(\FIFO[108][23] ), .IN3(\FIFO[110][23] ), .IN2(
        \FIFO[109][23] ), .IN4(\FIFO[111][23] ), .S0(n5850), .S1(n5944), .Q(
        n5350) );
  MUX41X1 U6324 ( .IN1(\FIFO[104][23] ), .IN3(\FIFO[106][23] ), .IN2(
        \FIFO[105][23] ), .IN4(\FIFO[107][23] ), .S0(n5850), .S1(n5944), .Q(
        n5351) );
  MUX41X1 U6325 ( .IN1(\FIFO[100][23] ), .IN3(\FIFO[102][23] ), .IN2(
        \FIFO[101][23] ), .IN4(\FIFO[103][23] ), .S0(n5850), .S1(n5944), .Q(
        n5352) );
  MUX41X1 U6326 ( .IN1(\FIFO[96][23] ), .IN3(\FIFO[98][23] ), .IN2(
        \FIFO[97][23] ), .IN4(\FIFO[99][23] ), .S0(n5850), .S1(n5944), .Q(
        n5353) );
  MUX41X1 U6327 ( .IN1(n5353), .IN3(n5351), .IN2(n5352), .IN4(n5350), .S0(
        n5750), .S1(n5769), .Q(n5354) );
  MUX41X1 U6328 ( .IN1(\FIFO[92][23] ), .IN3(\FIFO[94][23] ), .IN2(
        \FIFO[93][23] ), .IN4(\FIFO[95][23] ), .S0(n5850), .S1(n5944), .Q(
        n5355) );
  MUX41X1 U6329 ( .IN1(\FIFO[88][23] ), .IN3(\FIFO[90][23] ), .IN2(
        \FIFO[89][23] ), .IN4(\FIFO[91][23] ), .S0(n5850), .S1(n5944), .Q(
        n5356) );
  MUX41X1 U6330 ( .IN1(\FIFO[84][23] ), .IN3(\FIFO[86][23] ), .IN2(
        \FIFO[85][23] ), .IN4(\FIFO[87][23] ), .S0(n5850), .S1(n5944), .Q(
        n5357) );
  MUX41X1 U6331 ( .IN1(\FIFO[80][23] ), .IN3(\FIFO[82][23] ), .IN2(
        \FIFO[81][23] ), .IN4(\FIFO[83][23] ), .S0(n5850), .S1(n5944), .Q(
        n5358) );
  MUX41X1 U6332 ( .IN1(n5358), .IN3(n5356), .IN2(n5357), .IN4(n5355), .S0(
        n5750), .S1(n5769), .Q(n5359) );
  MUX41X1 U6333 ( .IN1(\FIFO[76][23] ), .IN3(\FIFO[78][23] ), .IN2(
        \FIFO[77][23] ), .IN4(\FIFO[79][23] ), .S0(n5851), .S1(n5945), .Q(
        n5360) );
  MUX41X1 U6334 ( .IN1(\FIFO[72][23] ), .IN3(\FIFO[74][23] ), .IN2(
        \FIFO[73][23] ), .IN4(\FIFO[75][23] ), .S0(n5851), .S1(n5945), .Q(
        n5361) );
  MUX41X1 U6335 ( .IN1(\FIFO[68][23] ), .IN3(\FIFO[70][23] ), .IN2(
        \FIFO[69][23] ), .IN4(\FIFO[71][23] ), .S0(n5851), .S1(n5945), .Q(
        n5362) );
  MUX41X1 U6336 ( .IN1(\FIFO[64][23] ), .IN3(\FIFO[66][23] ), .IN2(
        \FIFO[65][23] ), .IN4(\FIFO[67][23] ), .S0(n5851), .S1(n5945), .Q(
        n5363) );
  MUX41X1 U6337 ( .IN1(n5363), .IN3(n5361), .IN2(n5362), .IN4(n5360), .S0(
        n5750), .S1(n5769), .Q(n5364) );
  MUX41X1 U6338 ( .IN1(n5364), .IN3(n5354), .IN2(n5359), .IN4(n5349), .S0(
        n5729), .S1(n5733), .Q(n5365) );
  MUX41X1 U6339 ( .IN1(\FIFO[60][23] ), .IN3(\FIFO[62][23] ), .IN2(
        \FIFO[61][23] ), .IN4(\FIFO[63][23] ), .S0(n5851), .S1(n5945), .Q(
        n5366) );
  MUX41X1 U6340 ( .IN1(\FIFO[56][23] ), .IN3(\FIFO[58][23] ), .IN2(
        \FIFO[57][23] ), .IN4(\FIFO[59][23] ), .S0(n5851), .S1(n5945), .Q(
        n5367) );
  MUX41X1 U6341 ( .IN1(\FIFO[52][23] ), .IN3(\FIFO[54][23] ), .IN2(
        \FIFO[53][23] ), .IN4(\FIFO[55][23] ), .S0(n5851), .S1(n5945), .Q(
        n5368) );
  MUX41X1 U6342 ( .IN1(\FIFO[48][23] ), .IN3(\FIFO[50][23] ), .IN2(
        \FIFO[49][23] ), .IN4(\FIFO[51][23] ), .S0(n5851), .S1(n5945), .Q(
        n5369) );
  MUX41X1 U6343 ( .IN1(n5369), .IN3(n5367), .IN2(n5368), .IN4(n5366), .S0(
        n5750), .S1(n5769), .Q(n5370) );
  MUX41X1 U6344 ( .IN1(\FIFO[44][23] ), .IN3(\FIFO[46][23] ), .IN2(
        \FIFO[45][23] ), .IN4(\FIFO[47][23] ), .S0(n5851), .S1(n5945), .Q(
        n5371) );
  MUX41X1 U6345 ( .IN1(\FIFO[40][23] ), .IN3(\FIFO[42][23] ), .IN2(
        \FIFO[41][23] ), .IN4(\FIFO[43][23] ), .S0(n5851), .S1(n5945), .Q(
        n5372) );
  MUX41X1 U6346 ( .IN1(\FIFO[36][23] ), .IN3(\FIFO[38][23] ), .IN2(
        \FIFO[37][23] ), .IN4(\FIFO[39][23] ), .S0(n5851), .S1(n5945), .Q(
        n5373) );
  MUX41X1 U6347 ( .IN1(\FIFO[32][23] ), .IN3(\FIFO[34][23] ), .IN2(
        \FIFO[33][23] ), .IN4(\FIFO[35][23] ), .S0(n5851), .S1(n5945), .Q(
        n5374) );
  MUX41X1 U6348 ( .IN1(n5374), .IN3(n5372), .IN2(n5373), .IN4(n5371), .S0(
        n5750), .S1(n5769), .Q(n5375) );
  MUX41X1 U6349 ( .IN1(\FIFO[28][23] ), .IN3(\FIFO[30][23] ), .IN2(
        \FIFO[29][23] ), .IN4(\FIFO[31][23] ), .S0(n5852), .S1(n5946), .Q(
        n5376) );
  MUX41X1 U6350 ( .IN1(\FIFO[24][23] ), .IN3(\FIFO[26][23] ), .IN2(
        \FIFO[25][23] ), .IN4(\FIFO[27][23] ), .S0(n5852), .S1(n5946), .Q(
        n5377) );
  MUX41X1 U6351 ( .IN1(\FIFO[20][23] ), .IN3(\FIFO[22][23] ), .IN2(
        \FIFO[21][23] ), .IN4(\FIFO[23][23] ), .S0(n5852), .S1(n5946), .Q(
        n5378) );
  MUX41X1 U6352 ( .IN1(\FIFO[16][23] ), .IN3(\FIFO[18][23] ), .IN2(
        \FIFO[17][23] ), .IN4(\FIFO[19][23] ), .S0(n5852), .S1(n5946), .Q(
        n5379) );
  MUX41X1 U6353 ( .IN1(n5379), .IN3(n5377), .IN2(n5378), .IN4(n5376), .S0(
        n5750), .S1(n5769), .Q(n5380) );
  MUX41X1 U6354 ( .IN1(\FIFO[12][23] ), .IN3(\FIFO[14][23] ), .IN2(
        \FIFO[13][23] ), .IN4(\FIFO[15][23] ), .S0(n5852), .S1(n5946), .Q(
        n5381) );
  MUX41X1 U6355 ( .IN1(\FIFO[8][23] ), .IN3(\FIFO[10][23] ), .IN2(
        \FIFO[9][23] ), .IN4(\FIFO[11][23] ), .S0(n5852), .S1(n5946), .Q(n5382) );
  MUX41X1 U6356 ( .IN1(\FIFO[4][23] ), .IN3(\FIFO[6][23] ), .IN2(\FIFO[5][23] ), .IN4(\FIFO[7][23] ), .S0(n5852), .S1(n5946), .Q(n5383) );
  MUX41X1 U6357 ( .IN1(\FIFO[0][23] ), .IN3(\FIFO[2][23] ), .IN2(\FIFO[1][23] ), .IN4(\FIFO[3][23] ), .S0(n5852), .S1(n5946), .Q(n5384) );
  MUX41X1 U6358 ( .IN1(n5384), .IN3(n5382), .IN2(n5383), .IN4(n5381), .S0(
        n5750), .S1(n5769), .Q(n5385) );
  MUX41X1 U6359 ( .IN1(n5385), .IN3(n5375), .IN2(n5380), .IN4(n5370), .S0(
        n5729), .S1(n5733), .Q(n5386) );
  MUX21X1 U6360 ( .IN1(n5386), .IN2(n5365), .S(n5724), .Q(N227) );
  MUX41X1 U6361 ( .IN1(\FIFO[124][24] ), .IN3(\FIFO[126][24] ), .IN2(
        \FIFO[125][24] ), .IN4(\FIFO[127][24] ), .S0(n5852), .S1(n5946), .Q(
        n5387) );
  MUX41X1 U6362 ( .IN1(\FIFO[120][24] ), .IN3(\FIFO[122][24] ), .IN2(
        \FIFO[121][24] ), .IN4(\FIFO[123][24] ), .S0(n5852), .S1(n5946), .Q(
        n5388) );
  MUX41X1 U6363 ( .IN1(\FIFO[116][24] ), .IN3(\FIFO[118][24] ), .IN2(
        \FIFO[117][24] ), .IN4(\FIFO[119][24] ), .S0(n5852), .S1(n5946), .Q(
        n5389) );
  MUX41X1 U6364 ( .IN1(\FIFO[112][24] ), .IN3(\FIFO[114][24] ), .IN2(
        \FIFO[113][24] ), .IN4(\FIFO[115][24] ), .S0(n5852), .S1(n5946), .Q(
        n5390) );
  MUX41X1 U6365 ( .IN1(n5390), .IN3(n5388), .IN2(n5389), .IN4(n5387), .S0(
        n5750), .S1(n5769), .Q(n5391) );
  MUX41X1 U6366 ( .IN1(\FIFO[108][24] ), .IN3(\FIFO[110][24] ), .IN2(
        \FIFO[109][24] ), .IN4(\FIFO[111][24] ), .S0(n5853), .S1(n5947), .Q(
        n5392) );
  MUX41X1 U6367 ( .IN1(\FIFO[104][24] ), .IN3(\FIFO[106][24] ), .IN2(
        \FIFO[105][24] ), .IN4(\FIFO[107][24] ), .S0(n5853), .S1(n5947), .Q(
        n5393) );
  MUX41X1 U6368 ( .IN1(\FIFO[100][24] ), .IN3(\FIFO[102][24] ), .IN2(
        \FIFO[101][24] ), .IN4(\FIFO[103][24] ), .S0(n5853), .S1(n5947), .Q(
        n5394) );
  MUX41X1 U6369 ( .IN1(\FIFO[96][24] ), .IN3(\FIFO[98][24] ), .IN2(
        \FIFO[97][24] ), .IN4(\FIFO[99][24] ), .S0(n5853), .S1(n5947), .Q(
        n5395) );
  MUX41X1 U6370 ( .IN1(n5395), .IN3(n5393), .IN2(n5394), .IN4(n5392), .S0(
        n5750), .S1(n5769), .Q(n5396) );
  MUX41X1 U6371 ( .IN1(\FIFO[92][24] ), .IN3(\FIFO[94][24] ), .IN2(
        \FIFO[93][24] ), .IN4(\FIFO[95][24] ), .S0(n5853), .S1(n5947), .Q(
        n5397) );
  MUX41X1 U6372 ( .IN1(\FIFO[88][24] ), .IN3(\FIFO[90][24] ), .IN2(
        \FIFO[89][24] ), .IN4(\FIFO[91][24] ), .S0(n5853), .S1(n5947), .Q(
        n5398) );
  MUX41X1 U6373 ( .IN1(\FIFO[84][24] ), .IN3(\FIFO[86][24] ), .IN2(
        \FIFO[85][24] ), .IN4(\FIFO[87][24] ), .S0(n5853), .S1(n5947), .Q(
        n5399) );
  MUX41X1 U6374 ( .IN1(\FIFO[80][24] ), .IN3(\FIFO[82][24] ), .IN2(
        \FIFO[81][24] ), .IN4(\FIFO[83][24] ), .S0(n5853), .S1(n5947), .Q(
        n5400) );
  MUX41X1 U6375 ( .IN1(n5400), .IN3(n5398), .IN2(n5399), .IN4(n5397), .S0(
        n5750), .S1(n5769), .Q(n5401) );
  MUX41X1 U6376 ( .IN1(\FIFO[76][24] ), .IN3(\FIFO[78][24] ), .IN2(
        \FIFO[77][24] ), .IN4(\FIFO[79][24] ), .S0(n5853), .S1(n5947), .Q(
        n5402) );
  MUX41X1 U6377 ( .IN1(\FIFO[72][24] ), .IN3(\FIFO[74][24] ), .IN2(
        \FIFO[73][24] ), .IN4(\FIFO[75][24] ), .S0(n5853), .S1(n5947), .Q(
        n5403) );
  MUX41X1 U6378 ( .IN1(\FIFO[68][24] ), .IN3(\FIFO[70][24] ), .IN2(
        \FIFO[69][24] ), .IN4(\FIFO[71][24] ), .S0(n5853), .S1(n5947), .Q(
        n5404) );
  MUX41X1 U6379 ( .IN1(\FIFO[64][24] ), .IN3(\FIFO[66][24] ), .IN2(
        \FIFO[65][24] ), .IN4(\FIFO[67][24] ), .S0(n5853), .S1(n5947), .Q(
        n5405) );
  MUX41X1 U6380 ( .IN1(n5405), .IN3(n5403), .IN2(n5404), .IN4(n5402), .S0(
        n5750), .S1(n5769), .Q(n5406) );
  MUX41X1 U6381 ( .IN1(n5406), .IN3(n5396), .IN2(n5401), .IN4(n5391), .S0(
        n5729), .S1(n5733), .Q(n5407) );
  MUX41X1 U6382 ( .IN1(\FIFO[60][24] ), .IN3(\FIFO[62][24] ), .IN2(
        \FIFO[61][24] ), .IN4(\FIFO[63][24] ), .S0(n5854), .S1(n5948), .Q(
        n5408) );
  MUX41X1 U6383 ( .IN1(\FIFO[56][24] ), .IN3(\FIFO[58][24] ), .IN2(
        \FIFO[57][24] ), .IN4(\FIFO[59][24] ), .S0(n5854), .S1(n5948), .Q(
        n5409) );
  MUX41X1 U6384 ( .IN1(\FIFO[52][24] ), .IN3(\FIFO[54][24] ), .IN2(
        \FIFO[53][24] ), .IN4(\FIFO[55][24] ), .S0(n5854), .S1(n5948), .Q(
        n5410) );
  MUX41X1 U6385 ( .IN1(\FIFO[48][24] ), .IN3(\FIFO[50][24] ), .IN2(
        \FIFO[49][24] ), .IN4(\FIFO[51][24] ), .S0(n5854), .S1(n5948), .Q(
        n5411) );
  MUX41X1 U6386 ( .IN1(n5411), .IN3(n5409), .IN2(n5410), .IN4(n5408), .S0(
        n5751), .S1(n5770), .Q(n5412) );
  MUX41X1 U6387 ( .IN1(\FIFO[44][24] ), .IN3(\FIFO[46][24] ), .IN2(
        \FIFO[45][24] ), .IN4(\FIFO[47][24] ), .S0(n5854), .S1(n5948), .Q(
        n5413) );
  MUX41X1 U6388 ( .IN1(\FIFO[40][24] ), .IN3(\FIFO[42][24] ), .IN2(
        \FIFO[41][24] ), .IN4(\FIFO[43][24] ), .S0(n5854), .S1(n5948), .Q(
        n5414) );
  MUX41X1 U6389 ( .IN1(\FIFO[36][24] ), .IN3(\FIFO[38][24] ), .IN2(
        \FIFO[37][24] ), .IN4(\FIFO[39][24] ), .S0(n5854), .S1(n5948), .Q(
        n5415) );
  MUX41X1 U6390 ( .IN1(\FIFO[32][24] ), .IN3(\FIFO[34][24] ), .IN2(
        \FIFO[33][24] ), .IN4(\FIFO[35][24] ), .S0(n5854), .S1(n5948), .Q(
        n5416) );
  MUX41X1 U6391 ( .IN1(n5416), .IN3(n5414), .IN2(n5415), .IN4(n5413), .S0(
        n5751), .S1(n5770), .Q(n5417) );
  MUX41X1 U6392 ( .IN1(\FIFO[28][24] ), .IN3(\FIFO[30][24] ), .IN2(
        \FIFO[29][24] ), .IN4(\FIFO[31][24] ), .S0(n5854), .S1(n5948), .Q(
        n5418) );
  MUX41X1 U6393 ( .IN1(\FIFO[24][24] ), .IN3(\FIFO[26][24] ), .IN2(
        \FIFO[25][24] ), .IN4(\FIFO[27][24] ), .S0(n5854), .S1(n5948), .Q(
        n5419) );
  MUX41X1 U6394 ( .IN1(\FIFO[20][24] ), .IN3(\FIFO[22][24] ), .IN2(
        \FIFO[21][24] ), .IN4(\FIFO[23][24] ), .S0(n5854), .S1(n5948), .Q(
        n5420) );
  MUX41X1 U6395 ( .IN1(\FIFO[16][24] ), .IN3(\FIFO[18][24] ), .IN2(
        \FIFO[17][24] ), .IN4(\FIFO[19][24] ), .S0(n5854), .S1(n5948), .Q(
        n5421) );
  MUX41X1 U6396 ( .IN1(n5421), .IN3(n5419), .IN2(n5420), .IN4(n5418), .S0(
        n5751), .S1(n5770), .Q(n5422) );
  MUX41X1 U6397 ( .IN1(\FIFO[12][24] ), .IN3(\FIFO[14][24] ), .IN2(
        \FIFO[13][24] ), .IN4(\FIFO[15][24] ), .S0(n5855), .S1(n5949), .Q(
        n5423) );
  MUX41X1 U6398 ( .IN1(\FIFO[8][24] ), .IN3(\FIFO[10][24] ), .IN2(
        \FIFO[9][24] ), .IN4(\FIFO[11][24] ), .S0(n5855), .S1(n5949), .Q(n5424) );
  MUX41X1 U6399 ( .IN1(\FIFO[4][24] ), .IN3(\FIFO[6][24] ), .IN2(\FIFO[5][24] ), .IN4(\FIFO[7][24] ), .S0(n5855), .S1(n5949), .Q(n5425) );
  MUX41X1 U6400 ( .IN1(\FIFO[0][24] ), .IN3(\FIFO[2][24] ), .IN2(\FIFO[1][24] ), .IN4(\FIFO[3][24] ), .S0(n5855), .S1(n5949), .Q(n5426) );
  MUX41X1 U6401 ( .IN1(n5426), .IN3(n5424), .IN2(n5425), .IN4(n5423), .S0(
        n5751), .S1(n5770), .Q(n5427) );
  MUX41X1 U6402 ( .IN1(n5427), .IN3(n5417), .IN2(n5422), .IN4(n5412), .S0(
        n5729), .S1(n5733), .Q(n5428) );
  MUX21X1 U6403 ( .IN1(n5428), .IN2(n5407), .S(n5724), .Q(N226) );
  MUX41X1 U6404 ( .IN1(\FIFO[124][25] ), .IN3(\FIFO[126][25] ), .IN2(
        \FIFO[125][25] ), .IN4(\FIFO[127][25] ), .S0(n5855), .S1(n5949), .Q(
        n5429) );
  MUX41X1 U6405 ( .IN1(\FIFO[120][25] ), .IN3(\FIFO[122][25] ), .IN2(
        \FIFO[121][25] ), .IN4(\FIFO[123][25] ), .S0(n5855), .S1(n5949), .Q(
        n5430) );
  MUX41X1 U6406 ( .IN1(\FIFO[116][25] ), .IN3(\FIFO[118][25] ), .IN2(
        \FIFO[117][25] ), .IN4(\FIFO[119][25] ), .S0(n5855), .S1(n5949), .Q(
        n5431) );
  MUX41X1 U6407 ( .IN1(\FIFO[112][25] ), .IN3(\FIFO[114][25] ), .IN2(
        \FIFO[113][25] ), .IN4(\FIFO[115][25] ), .S0(n5855), .S1(n5949), .Q(
        n5432) );
  MUX41X1 U6408 ( .IN1(n5432), .IN3(n5430), .IN2(n5431), .IN4(n5429), .S0(
        n5751), .S1(n5770), .Q(n5433) );
  MUX41X1 U6409 ( .IN1(\FIFO[108][25] ), .IN3(\FIFO[110][25] ), .IN2(
        \FIFO[109][25] ), .IN4(\FIFO[111][25] ), .S0(n5855), .S1(n5949), .Q(
        n5434) );
  MUX41X1 U6410 ( .IN1(\FIFO[104][25] ), .IN3(\FIFO[106][25] ), .IN2(
        \FIFO[105][25] ), .IN4(\FIFO[107][25] ), .S0(n5855), .S1(n5949), .Q(
        n5435) );
  MUX41X1 U6411 ( .IN1(\FIFO[100][25] ), .IN3(\FIFO[102][25] ), .IN2(
        \FIFO[101][25] ), .IN4(\FIFO[103][25] ), .S0(n5855), .S1(n5949), .Q(
        n5436) );
  MUX41X1 U6412 ( .IN1(\FIFO[96][25] ), .IN3(\FIFO[98][25] ), .IN2(
        \FIFO[97][25] ), .IN4(\FIFO[99][25] ), .S0(n5855), .S1(n5949), .Q(
        n5437) );
  MUX41X1 U6413 ( .IN1(n5437), .IN3(n5435), .IN2(n5436), .IN4(n5434), .S0(
        n5751), .S1(n5770), .Q(n5438) );
  MUX41X1 U6414 ( .IN1(\FIFO[92][25] ), .IN3(\FIFO[94][25] ), .IN2(
        \FIFO[93][25] ), .IN4(\FIFO[95][25] ), .S0(n5856), .S1(n5950), .Q(
        n5439) );
  MUX41X1 U6415 ( .IN1(\FIFO[88][25] ), .IN3(\FIFO[90][25] ), .IN2(
        \FIFO[89][25] ), .IN4(\FIFO[91][25] ), .S0(n5856), .S1(n5950), .Q(
        n5440) );
  MUX41X1 U6416 ( .IN1(\FIFO[84][25] ), .IN3(\FIFO[86][25] ), .IN2(
        \FIFO[85][25] ), .IN4(\FIFO[87][25] ), .S0(n5856), .S1(n5950), .Q(
        n5441) );
  MUX41X1 U6417 ( .IN1(\FIFO[80][25] ), .IN3(\FIFO[82][25] ), .IN2(
        \FIFO[81][25] ), .IN4(\FIFO[83][25] ), .S0(n5856), .S1(n5950), .Q(
        n5442) );
  MUX41X1 U6418 ( .IN1(n5442), .IN3(n5440), .IN2(n5441), .IN4(n5439), .S0(
        n5751), .S1(n5770), .Q(n5443) );
  MUX41X1 U6419 ( .IN1(\FIFO[76][25] ), .IN3(\FIFO[78][25] ), .IN2(
        \FIFO[77][25] ), .IN4(\FIFO[79][25] ), .S0(n5856), .S1(n5950), .Q(
        n5444) );
  MUX41X1 U6420 ( .IN1(\FIFO[72][25] ), .IN3(\FIFO[74][25] ), .IN2(
        \FIFO[73][25] ), .IN4(\FIFO[75][25] ), .S0(n5856), .S1(n5950), .Q(
        n5445) );
  MUX41X1 U6421 ( .IN1(\FIFO[68][25] ), .IN3(\FIFO[70][25] ), .IN2(
        \FIFO[69][25] ), .IN4(\FIFO[71][25] ), .S0(n5856), .S1(n5950), .Q(
        n5446) );
  MUX41X1 U6422 ( .IN1(\FIFO[64][25] ), .IN3(\FIFO[66][25] ), .IN2(
        \FIFO[65][25] ), .IN4(\FIFO[67][25] ), .S0(n5856), .S1(n5950), .Q(
        n5447) );
  MUX41X1 U6423 ( .IN1(n5447), .IN3(n5445), .IN2(n5446), .IN4(n5444), .S0(
        n5751), .S1(n5770), .Q(n5448) );
  MUX41X1 U6424 ( .IN1(n5448), .IN3(n5438), .IN2(n5443), .IN4(n5433), .S0(
        n5729), .S1(n5733), .Q(n5449) );
  MUX41X1 U6425 ( .IN1(\FIFO[60][25] ), .IN3(\FIFO[62][25] ), .IN2(
        \FIFO[61][25] ), .IN4(\FIFO[63][25] ), .S0(n5856), .S1(n5950), .Q(
        n5450) );
  MUX41X1 U6426 ( .IN1(\FIFO[56][25] ), .IN3(\FIFO[58][25] ), .IN2(
        \FIFO[57][25] ), .IN4(\FIFO[59][25] ), .S0(n5856), .S1(n5950), .Q(
        n5451) );
  MUX41X1 U6427 ( .IN1(\FIFO[52][25] ), .IN3(\FIFO[54][25] ), .IN2(
        \FIFO[53][25] ), .IN4(\FIFO[55][25] ), .S0(n5856), .S1(n5950), .Q(
        n5452) );
  MUX41X1 U6428 ( .IN1(\FIFO[48][25] ), .IN3(\FIFO[50][25] ), .IN2(
        \FIFO[49][25] ), .IN4(\FIFO[51][25] ), .S0(n5856), .S1(n5950), .Q(
        n5453) );
  MUX41X1 U6429 ( .IN1(n5453), .IN3(n5451), .IN2(n5452), .IN4(n5450), .S0(
        n5751), .S1(n5770), .Q(n5454) );
  MUX41X1 U6430 ( .IN1(\FIFO[44][25] ), .IN3(\FIFO[46][25] ), .IN2(
        \FIFO[45][25] ), .IN4(\FIFO[47][25] ), .S0(n5857), .S1(n5951), .Q(
        n5455) );
  MUX41X1 U6431 ( .IN1(\FIFO[40][25] ), .IN3(\FIFO[42][25] ), .IN2(
        \FIFO[41][25] ), .IN4(\FIFO[43][25] ), .S0(n5857), .S1(n5951), .Q(
        n5456) );
  MUX41X1 U6432 ( .IN1(\FIFO[36][25] ), .IN3(\FIFO[38][25] ), .IN2(
        \FIFO[37][25] ), .IN4(\FIFO[39][25] ), .S0(n5857), .S1(n5951), .Q(
        n5457) );
  MUX41X1 U6433 ( .IN1(\FIFO[32][25] ), .IN3(\FIFO[34][25] ), .IN2(
        \FIFO[33][25] ), .IN4(\FIFO[35][25] ), .S0(n5857), .S1(n5951), .Q(
        n5458) );
  MUX41X1 U6434 ( .IN1(n5458), .IN3(n5456), .IN2(n5457), .IN4(n5455), .S0(
        n5751), .S1(n5770), .Q(n5459) );
  MUX41X1 U6435 ( .IN1(\FIFO[28][25] ), .IN3(\FIFO[30][25] ), .IN2(
        \FIFO[29][25] ), .IN4(\FIFO[31][25] ), .S0(n5857), .S1(n5951), .Q(
        n5460) );
  MUX41X1 U6436 ( .IN1(\FIFO[24][25] ), .IN3(\FIFO[26][25] ), .IN2(
        \FIFO[25][25] ), .IN4(\FIFO[27][25] ), .S0(n5857), .S1(n5951), .Q(
        n5461) );
  MUX41X1 U6437 ( .IN1(\FIFO[20][25] ), .IN3(\FIFO[22][25] ), .IN2(
        \FIFO[21][25] ), .IN4(\FIFO[23][25] ), .S0(n5857), .S1(n5951), .Q(
        n5462) );
  MUX41X1 U6438 ( .IN1(\FIFO[16][25] ), .IN3(\FIFO[18][25] ), .IN2(
        \FIFO[17][25] ), .IN4(\FIFO[19][25] ), .S0(n5857), .S1(n5951), .Q(
        n5463) );
  MUX41X1 U6439 ( .IN1(n5463), .IN3(n5461), .IN2(n5462), .IN4(n5460), .S0(
        n5751), .S1(n5770), .Q(n5464) );
  MUX41X1 U6440 ( .IN1(\FIFO[12][25] ), .IN3(\FIFO[14][25] ), .IN2(
        \FIFO[13][25] ), .IN4(\FIFO[15][25] ), .S0(n5857), .S1(n5951), .Q(
        n5465) );
  MUX41X1 U6441 ( .IN1(\FIFO[8][25] ), .IN3(\FIFO[10][25] ), .IN2(
        \FIFO[9][25] ), .IN4(\FIFO[11][25] ), .S0(n5857), .S1(n5951), .Q(n5466) );
  MUX41X1 U6442 ( .IN1(\FIFO[4][25] ), .IN3(\FIFO[6][25] ), .IN2(\FIFO[5][25] ), .IN4(\FIFO[7][25] ), .S0(n5857), .S1(n5951), .Q(n5467) );
  MUX41X1 U6443 ( .IN1(\FIFO[0][25] ), .IN3(\FIFO[2][25] ), .IN2(\FIFO[1][25] ), .IN4(\FIFO[3][25] ), .S0(n5857), .S1(n5951), .Q(n5468) );
  MUX41X1 U6444 ( .IN1(n5468), .IN3(n5466), .IN2(n5467), .IN4(n5465), .S0(
        n5751), .S1(n5770), .Q(n5469) );
  MUX41X1 U6445 ( .IN1(n5469), .IN3(n5459), .IN2(n5464), .IN4(n5454), .S0(
        n5729), .S1(n5733), .Q(n5470) );
  MUX21X1 U6446 ( .IN1(n5470), .IN2(n5449), .S(n5724), .Q(N225) );
  MUX41X1 U6447 ( .IN1(\FIFO[124][26] ), .IN3(\FIFO[126][26] ), .IN2(
        \FIFO[125][26] ), .IN4(\FIFO[127][26] ), .S0(n5858), .S1(n5952), .Q(
        n5471) );
  MUX41X1 U6448 ( .IN1(\FIFO[120][26] ), .IN3(\FIFO[122][26] ), .IN2(
        \FIFO[121][26] ), .IN4(\FIFO[123][26] ), .S0(n5858), .S1(n5952), .Q(
        n5472) );
  MUX41X1 U6449 ( .IN1(\FIFO[116][26] ), .IN3(\FIFO[118][26] ), .IN2(
        \FIFO[117][26] ), .IN4(\FIFO[119][26] ), .S0(n5858), .S1(n5952), .Q(
        n5473) );
  MUX41X1 U6450 ( .IN1(\FIFO[112][26] ), .IN3(\FIFO[114][26] ), .IN2(
        \FIFO[113][26] ), .IN4(\FIFO[115][26] ), .S0(n5858), .S1(n5952), .Q(
        n5474) );
  MUX41X1 U6451 ( .IN1(n5474), .IN3(n5472), .IN2(n5473), .IN4(n5471), .S0(
        n5752), .S1(n5771), .Q(n5475) );
  MUX41X1 U6452 ( .IN1(\FIFO[108][26] ), .IN3(\FIFO[110][26] ), .IN2(
        \FIFO[109][26] ), .IN4(\FIFO[111][26] ), .S0(n5858), .S1(n5952), .Q(
        n5476) );
  MUX41X1 U6453 ( .IN1(\FIFO[104][26] ), .IN3(\FIFO[106][26] ), .IN2(
        \FIFO[105][26] ), .IN4(\FIFO[107][26] ), .S0(n5858), .S1(n5952), .Q(
        n5477) );
  MUX41X1 U6454 ( .IN1(\FIFO[100][26] ), .IN3(\FIFO[102][26] ), .IN2(
        \FIFO[101][26] ), .IN4(\FIFO[103][26] ), .S0(n5858), .S1(n5952), .Q(
        n5478) );
  MUX41X1 U6455 ( .IN1(\FIFO[96][26] ), .IN3(\FIFO[98][26] ), .IN2(
        \FIFO[97][26] ), .IN4(\FIFO[99][26] ), .S0(n5858), .S1(n5952), .Q(
        n5479) );
  MUX41X1 U6456 ( .IN1(n5479), .IN3(n5477), .IN2(n5478), .IN4(n5476), .S0(
        n5752), .S1(n5771), .Q(n5480) );
  MUX41X1 U6457 ( .IN1(\FIFO[92][26] ), .IN3(\FIFO[94][26] ), .IN2(
        \FIFO[93][26] ), .IN4(\FIFO[95][26] ), .S0(n5858), .S1(n5952), .Q(
        n5481) );
  MUX41X1 U6458 ( .IN1(\FIFO[88][26] ), .IN3(\FIFO[90][26] ), .IN2(
        \FIFO[89][26] ), .IN4(\FIFO[91][26] ), .S0(n5858), .S1(n5952), .Q(
        n5482) );
  MUX41X1 U6459 ( .IN1(\FIFO[84][26] ), .IN3(\FIFO[86][26] ), .IN2(
        \FIFO[85][26] ), .IN4(\FIFO[87][26] ), .S0(n5858), .S1(n5952), .Q(
        n5483) );
  MUX41X1 U6460 ( .IN1(\FIFO[80][26] ), .IN3(\FIFO[82][26] ), .IN2(
        \FIFO[81][26] ), .IN4(\FIFO[83][26] ), .S0(n5858), .S1(n5952), .Q(
        n5484) );
  MUX41X1 U6461 ( .IN1(n5484), .IN3(n5482), .IN2(n5483), .IN4(n5481), .S0(
        n5752), .S1(n5771), .Q(n5485) );
  MUX41X1 U6462 ( .IN1(\FIFO[76][26] ), .IN3(\FIFO[78][26] ), .IN2(
        \FIFO[77][26] ), .IN4(\FIFO[79][26] ), .S0(n5859), .S1(n5953), .Q(
        n5486) );
  MUX41X1 U6463 ( .IN1(\FIFO[72][26] ), .IN3(\FIFO[74][26] ), .IN2(
        \FIFO[73][26] ), .IN4(\FIFO[75][26] ), .S0(n5859), .S1(n5953), .Q(
        n5487) );
  MUX41X1 U6464 ( .IN1(\FIFO[68][26] ), .IN3(\FIFO[70][26] ), .IN2(
        \FIFO[69][26] ), .IN4(\FIFO[71][26] ), .S0(n5859), .S1(n5953), .Q(
        n5488) );
  MUX41X1 U6465 ( .IN1(\FIFO[64][26] ), .IN3(\FIFO[66][26] ), .IN2(
        \FIFO[65][26] ), .IN4(\FIFO[67][26] ), .S0(n5859), .S1(n5953), .Q(
        n5489) );
  MUX41X1 U6466 ( .IN1(n5489), .IN3(n5487), .IN2(n5488), .IN4(n5486), .S0(
        n5752), .S1(n5771), .Q(n5490) );
  MUX41X1 U6467 ( .IN1(n5490), .IN3(n5480), .IN2(n5485), .IN4(n5475), .S0(
        n5725), .S1(n5734), .Q(n5491) );
  MUX41X1 U6468 ( .IN1(\FIFO[60][26] ), .IN3(\FIFO[62][26] ), .IN2(
        \FIFO[61][26] ), .IN4(\FIFO[63][26] ), .S0(n5859), .S1(n5953), .Q(
        n5492) );
  MUX41X1 U6469 ( .IN1(\FIFO[56][26] ), .IN3(\FIFO[58][26] ), .IN2(
        \FIFO[57][26] ), .IN4(\FIFO[59][26] ), .S0(n5859), .S1(n5953), .Q(
        n5493) );
  MUX41X1 U6470 ( .IN1(\FIFO[52][26] ), .IN3(\FIFO[54][26] ), .IN2(
        \FIFO[53][26] ), .IN4(\FIFO[55][26] ), .S0(n5859), .S1(n5953), .Q(
        n5494) );
  MUX41X1 U6471 ( .IN1(\FIFO[48][26] ), .IN3(\FIFO[50][26] ), .IN2(
        \FIFO[49][26] ), .IN4(\FIFO[51][26] ), .S0(n5859), .S1(n5953), .Q(
        n5495) );
  MUX41X1 U6472 ( .IN1(n5495), .IN3(n5493), .IN2(n5494), .IN4(n5492), .S0(
        n5752), .S1(n5771), .Q(n5496) );
  MUX41X1 U6473 ( .IN1(\FIFO[44][26] ), .IN3(\FIFO[46][26] ), .IN2(
        \FIFO[45][26] ), .IN4(\FIFO[47][26] ), .S0(n5859), .S1(n5953), .Q(
        n5497) );
  MUX41X1 U6474 ( .IN1(\FIFO[40][26] ), .IN3(\FIFO[42][26] ), .IN2(
        \FIFO[41][26] ), .IN4(\FIFO[43][26] ), .S0(n5859), .S1(n5953), .Q(
        n5498) );
  MUX41X1 U6475 ( .IN1(\FIFO[36][26] ), .IN3(\FIFO[38][26] ), .IN2(
        \FIFO[37][26] ), .IN4(\FIFO[39][26] ), .S0(n5859), .S1(n5953), .Q(
        n5499) );
  MUX41X1 U6476 ( .IN1(\FIFO[32][26] ), .IN3(\FIFO[34][26] ), .IN2(
        \FIFO[33][26] ), .IN4(\FIFO[35][26] ), .S0(n5859), .S1(n5953), .Q(
        n5500) );
  MUX41X1 U6477 ( .IN1(n5500), .IN3(n5498), .IN2(n5499), .IN4(n5497), .S0(
        n5752), .S1(n5771), .Q(n5501) );
  MUX41X1 U6478 ( .IN1(\FIFO[28][26] ), .IN3(\FIFO[30][26] ), .IN2(
        \FIFO[29][26] ), .IN4(\FIFO[31][26] ), .S0(n5860), .S1(n5954), .Q(
        n5502) );
  MUX41X1 U6479 ( .IN1(\FIFO[24][26] ), .IN3(\FIFO[26][26] ), .IN2(
        \FIFO[25][26] ), .IN4(\FIFO[27][26] ), .S0(n5860), .S1(n5954), .Q(
        n5503) );
  MUX41X1 U6480 ( .IN1(\FIFO[20][26] ), .IN3(\FIFO[22][26] ), .IN2(
        \FIFO[21][26] ), .IN4(\FIFO[23][26] ), .S0(n5860), .S1(n5954), .Q(
        n5504) );
  MUX41X1 U6481 ( .IN1(\FIFO[16][26] ), .IN3(\FIFO[18][26] ), .IN2(
        \FIFO[17][26] ), .IN4(\FIFO[19][26] ), .S0(n5860), .S1(n5954), .Q(
        n5505) );
  MUX41X1 U6482 ( .IN1(n5505), .IN3(n5503), .IN2(n5504), .IN4(n5502), .S0(
        n5752), .S1(n5771), .Q(n5506) );
  MUX41X1 U6483 ( .IN1(\FIFO[12][26] ), .IN3(\FIFO[14][26] ), .IN2(
        \FIFO[13][26] ), .IN4(\FIFO[15][26] ), .S0(n5860), .S1(n5954), .Q(
        n5507) );
  MUX41X1 U6484 ( .IN1(\FIFO[8][26] ), .IN3(\FIFO[10][26] ), .IN2(
        \FIFO[9][26] ), .IN4(\FIFO[11][26] ), .S0(n5860), .S1(n5954), .Q(n5508) );
  MUX41X1 U6485 ( .IN1(\FIFO[4][26] ), .IN3(\FIFO[6][26] ), .IN2(\FIFO[5][26] ), .IN4(\FIFO[7][26] ), .S0(n5860), .S1(n5954), .Q(n5509) );
  MUX41X1 U6486 ( .IN1(\FIFO[0][26] ), .IN3(\FIFO[2][26] ), .IN2(\FIFO[1][26] ), .IN4(\FIFO[3][26] ), .S0(n5860), .S1(n5954), .Q(n5510) );
  MUX41X1 U6487 ( .IN1(n5510), .IN3(n5508), .IN2(n5509), .IN4(n5507), .S0(
        n5752), .S1(n5771), .Q(n5511) );
  MUX41X1 U6488 ( .IN1(n5511), .IN3(n5501), .IN2(n5506), .IN4(n5496), .S0(
        n5725), .S1(n5734), .Q(n5512) );
  MUX21X1 U6489 ( .IN1(n5512), .IN2(n5491), .S(n5724), .Q(N224) );
  MUX41X1 U6490 ( .IN1(\FIFO[124][27] ), .IN3(\FIFO[126][27] ), .IN2(
        \FIFO[125][27] ), .IN4(\FIFO[127][27] ), .S0(n5860), .S1(n5954), .Q(
        n5513) );
  MUX41X1 U6491 ( .IN1(\FIFO[120][27] ), .IN3(\FIFO[122][27] ), .IN2(
        \FIFO[121][27] ), .IN4(\FIFO[123][27] ), .S0(n5860), .S1(n5954), .Q(
        n5514) );
  MUX41X1 U6492 ( .IN1(\FIFO[116][27] ), .IN3(\FIFO[118][27] ), .IN2(
        \FIFO[117][27] ), .IN4(\FIFO[119][27] ), .S0(n5860), .S1(n5954), .Q(
        n5515) );
  MUX41X1 U6493 ( .IN1(\FIFO[112][27] ), .IN3(\FIFO[114][27] ), .IN2(
        \FIFO[113][27] ), .IN4(\FIFO[115][27] ), .S0(n5860), .S1(n5954), .Q(
        n5516) );
  MUX41X1 U6494 ( .IN1(n5516), .IN3(n5514), .IN2(n5515), .IN4(n5513), .S0(
        n5752), .S1(n5771), .Q(n5517) );
  MUX41X1 U6495 ( .IN1(\FIFO[108][27] ), .IN3(\FIFO[110][27] ), .IN2(
        \FIFO[109][27] ), .IN4(\FIFO[111][27] ), .S0(n5861), .S1(n5955), .Q(
        n5518) );
  MUX41X1 U6496 ( .IN1(\FIFO[104][27] ), .IN3(\FIFO[106][27] ), .IN2(
        \FIFO[105][27] ), .IN4(\FIFO[107][27] ), .S0(n5861), .S1(n5955), .Q(
        n5519) );
  MUX41X1 U6497 ( .IN1(\FIFO[100][27] ), .IN3(\FIFO[102][27] ), .IN2(
        \FIFO[101][27] ), .IN4(\FIFO[103][27] ), .S0(n5861), .S1(n5955), .Q(
        n5520) );
  MUX41X1 U6498 ( .IN1(\FIFO[96][27] ), .IN3(\FIFO[98][27] ), .IN2(
        \FIFO[97][27] ), .IN4(\FIFO[99][27] ), .S0(n5861), .S1(n5955), .Q(
        n5521) );
  MUX41X1 U6499 ( .IN1(n5521), .IN3(n5519), .IN2(n5520), .IN4(n5518), .S0(
        n5752), .S1(n5771), .Q(n5522) );
  MUX41X1 U6500 ( .IN1(\FIFO[92][27] ), .IN3(\FIFO[94][27] ), .IN2(
        \FIFO[93][27] ), .IN4(\FIFO[95][27] ), .S0(n5861), .S1(n5955), .Q(
        n5523) );
  MUX41X1 U6501 ( .IN1(\FIFO[88][27] ), .IN3(\FIFO[90][27] ), .IN2(
        \FIFO[89][27] ), .IN4(\FIFO[91][27] ), .S0(n5861), .S1(n5955), .Q(
        n5524) );
  MUX41X1 U6502 ( .IN1(\FIFO[84][27] ), .IN3(\FIFO[86][27] ), .IN2(
        \FIFO[85][27] ), .IN4(\FIFO[87][27] ), .S0(n5861), .S1(n5955), .Q(
        n5525) );
  MUX41X1 U6503 ( .IN1(\FIFO[80][27] ), .IN3(\FIFO[82][27] ), .IN2(
        \FIFO[81][27] ), .IN4(\FIFO[83][27] ), .S0(n5861), .S1(n5955), .Q(
        n5526) );
  MUX41X1 U6504 ( .IN1(n5526), .IN3(n5524), .IN2(n5525), .IN4(n5523), .S0(
        n5752), .S1(n5771), .Q(n5527) );
  MUX41X1 U6505 ( .IN1(\FIFO[76][27] ), .IN3(\FIFO[78][27] ), .IN2(
        \FIFO[77][27] ), .IN4(\FIFO[79][27] ), .S0(n5861), .S1(n5955), .Q(
        n5528) );
  MUX41X1 U6506 ( .IN1(\FIFO[72][27] ), .IN3(\FIFO[74][27] ), .IN2(
        \FIFO[73][27] ), .IN4(\FIFO[75][27] ), .S0(n5861), .S1(n5955), .Q(
        n5529) );
  MUX41X1 U6507 ( .IN1(\FIFO[68][27] ), .IN3(\FIFO[70][27] ), .IN2(
        \FIFO[69][27] ), .IN4(\FIFO[71][27] ), .S0(n5861), .S1(n5955), .Q(
        n5530) );
  MUX41X1 U6508 ( .IN1(\FIFO[64][27] ), .IN3(\FIFO[66][27] ), .IN2(
        \FIFO[65][27] ), .IN4(\FIFO[67][27] ), .S0(n5861), .S1(n5955), .Q(
        n5531) );
  MUX41X1 U6509 ( .IN1(n5531), .IN3(n5529), .IN2(n5530), .IN4(n5528), .S0(
        n5752), .S1(n5771), .Q(n5532) );
  MUX41X1 U6510 ( .IN1(n5532), .IN3(n5522), .IN2(n5527), .IN4(n5517), .S0(
        n5725), .S1(n5734), .Q(n5533) );
  MUX41X1 U6511 ( .IN1(\FIFO[60][27] ), .IN3(\FIFO[62][27] ), .IN2(
        \FIFO[61][27] ), .IN4(\FIFO[63][27] ), .S0(n5862), .S1(n5956), .Q(
        n5534) );
  MUX41X1 U6512 ( .IN1(\FIFO[56][27] ), .IN3(\FIFO[58][27] ), .IN2(
        \FIFO[57][27] ), .IN4(\FIFO[59][27] ), .S0(n5862), .S1(n5956), .Q(
        n5535) );
  MUX41X1 U6513 ( .IN1(\FIFO[52][27] ), .IN3(\FIFO[54][27] ), .IN2(
        \FIFO[53][27] ), .IN4(\FIFO[55][27] ), .S0(n5862), .S1(n5956), .Q(
        n5536) );
  MUX41X1 U6514 ( .IN1(\FIFO[48][27] ), .IN3(\FIFO[50][27] ), .IN2(
        \FIFO[49][27] ), .IN4(\FIFO[51][27] ), .S0(n5862), .S1(n5956), .Q(
        n5537) );
  MUX41X1 U6515 ( .IN1(n5537), .IN3(n5535), .IN2(n5536), .IN4(n5534), .S0(
        n5753), .S1(n5772), .Q(n5538) );
  MUX41X1 U6516 ( .IN1(\FIFO[44][27] ), .IN3(\FIFO[46][27] ), .IN2(
        \FIFO[45][27] ), .IN4(\FIFO[47][27] ), .S0(n5862), .S1(n5956), .Q(
        n5539) );
  MUX41X1 U6517 ( .IN1(\FIFO[40][27] ), .IN3(\FIFO[42][27] ), .IN2(
        \FIFO[41][27] ), .IN4(\FIFO[43][27] ), .S0(n5862), .S1(n5956), .Q(
        n5540) );
  MUX41X1 U6518 ( .IN1(\FIFO[36][27] ), .IN3(\FIFO[38][27] ), .IN2(
        \FIFO[37][27] ), .IN4(\FIFO[39][27] ), .S0(n5862), .S1(n5956), .Q(
        n5541) );
  MUX41X1 U6519 ( .IN1(\FIFO[32][27] ), .IN3(\FIFO[34][27] ), .IN2(
        \FIFO[33][27] ), .IN4(\FIFO[35][27] ), .S0(n5862), .S1(n5956), .Q(
        n5542) );
  MUX41X1 U6520 ( .IN1(n5542), .IN3(n5540), .IN2(n5541), .IN4(n5539), .S0(
        n5753), .S1(n5772), .Q(n5543) );
  MUX41X1 U6521 ( .IN1(\FIFO[28][27] ), .IN3(\FIFO[30][27] ), .IN2(
        \FIFO[29][27] ), .IN4(\FIFO[31][27] ), .S0(n5862), .S1(n5956), .Q(
        n5544) );
  MUX41X1 U6522 ( .IN1(\FIFO[24][27] ), .IN3(\FIFO[26][27] ), .IN2(
        \FIFO[25][27] ), .IN4(\FIFO[27][27] ), .S0(n5862), .S1(n5956), .Q(
        n5545) );
  MUX41X1 U6523 ( .IN1(\FIFO[20][27] ), .IN3(\FIFO[22][27] ), .IN2(
        \FIFO[21][27] ), .IN4(\FIFO[23][27] ), .S0(n5862), .S1(n5956), .Q(
        n5546) );
  MUX41X1 U6524 ( .IN1(\FIFO[16][27] ), .IN3(\FIFO[18][27] ), .IN2(
        \FIFO[17][27] ), .IN4(\FIFO[19][27] ), .S0(n5862), .S1(n5956), .Q(
        n5547) );
  MUX41X1 U6525 ( .IN1(n5547), .IN3(n5545), .IN2(n5546), .IN4(n5544), .S0(
        n5753), .S1(n5772), .Q(n5548) );
  MUX41X1 U6526 ( .IN1(\FIFO[12][27] ), .IN3(\FIFO[14][27] ), .IN2(
        \FIFO[13][27] ), .IN4(\FIFO[15][27] ), .S0(n5863), .S1(n5957), .Q(
        n5549) );
  MUX41X1 U6527 ( .IN1(\FIFO[8][27] ), .IN3(\FIFO[10][27] ), .IN2(
        \FIFO[9][27] ), .IN4(\FIFO[11][27] ), .S0(n5863), .S1(n5957), .Q(n5550) );
  MUX41X1 U6528 ( .IN1(\FIFO[4][27] ), .IN3(\FIFO[6][27] ), .IN2(\FIFO[5][27] ), .IN4(\FIFO[7][27] ), .S0(n5863), .S1(n5957), .Q(n5551) );
  MUX41X1 U6529 ( .IN1(\FIFO[0][27] ), .IN3(\FIFO[2][27] ), .IN2(\FIFO[1][27] ), .IN4(\FIFO[3][27] ), .S0(n5863), .S1(n5957), .Q(n5552) );
  MUX41X1 U6530 ( .IN1(n5552), .IN3(n5550), .IN2(n5551), .IN4(n5549), .S0(
        n5753), .S1(n5772), .Q(n5553) );
  MUX41X1 U6531 ( .IN1(n5553), .IN3(n5543), .IN2(n5548), .IN4(n5538), .S0(
        n5726), .S1(n5734), .Q(n5554) );
  MUX21X1 U6532 ( .IN1(n5554), .IN2(n5533), .S(n5724), .Q(N223) );
  MUX41X1 U6533 ( .IN1(\FIFO[124][28] ), .IN3(\FIFO[126][28] ), .IN2(
        \FIFO[125][28] ), .IN4(\FIFO[127][28] ), .S0(n5863), .S1(n5957), .Q(
        n5555) );
  MUX41X1 U6534 ( .IN1(\FIFO[120][28] ), .IN3(\FIFO[122][28] ), .IN2(
        \FIFO[121][28] ), .IN4(\FIFO[123][28] ), .S0(n5863), .S1(n5957), .Q(
        n5556) );
  MUX41X1 U6535 ( .IN1(\FIFO[116][28] ), .IN3(\FIFO[118][28] ), .IN2(
        \FIFO[117][28] ), .IN4(\FIFO[119][28] ), .S0(n5863), .S1(n5957), .Q(
        n5557) );
  MUX41X1 U6536 ( .IN1(\FIFO[112][28] ), .IN3(\FIFO[114][28] ), .IN2(
        \FIFO[113][28] ), .IN4(\FIFO[115][28] ), .S0(n5863), .S1(n5957), .Q(
        n5558) );
  MUX41X1 U6537 ( .IN1(n5558), .IN3(n5556), .IN2(n5557), .IN4(n5555), .S0(
        n5753), .S1(n5772), .Q(n5559) );
  MUX41X1 U6538 ( .IN1(\FIFO[108][28] ), .IN3(\FIFO[110][28] ), .IN2(
        \FIFO[109][28] ), .IN4(\FIFO[111][28] ), .S0(n5863), .S1(n5957), .Q(
        n5560) );
  MUX41X1 U6539 ( .IN1(\FIFO[104][28] ), .IN3(\FIFO[106][28] ), .IN2(
        \FIFO[105][28] ), .IN4(\FIFO[107][28] ), .S0(n5863), .S1(n5957), .Q(
        n5561) );
  MUX41X1 U6540 ( .IN1(\FIFO[100][28] ), .IN3(\FIFO[102][28] ), .IN2(
        \FIFO[101][28] ), .IN4(\FIFO[103][28] ), .S0(n5863), .S1(n5957), .Q(
        n5562) );
  MUX41X1 U6541 ( .IN1(\FIFO[96][28] ), .IN3(\FIFO[98][28] ), .IN2(
        \FIFO[97][28] ), .IN4(\FIFO[99][28] ), .S0(n5863), .S1(n5957), .Q(
        n5563) );
  MUX41X1 U6542 ( .IN1(n5563), .IN3(n5561), .IN2(n5562), .IN4(n5560), .S0(
        n5753), .S1(n5772), .Q(n5564) );
  MUX41X1 U6543 ( .IN1(\FIFO[92][28] ), .IN3(\FIFO[94][28] ), .IN2(
        \FIFO[93][28] ), .IN4(\FIFO[95][28] ), .S0(n5864), .S1(n5958), .Q(
        n5565) );
  MUX41X1 U6544 ( .IN1(\FIFO[88][28] ), .IN3(\FIFO[90][28] ), .IN2(
        \FIFO[89][28] ), .IN4(\FIFO[91][28] ), .S0(n5864), .S1(n5958), .Q(
        n5566) );
  MUX41X1 U6545 ( .IN1(\FIFO[84][28] ), .IN3(\FIFO[86][28] ), .IN2(
        \FIFO[85][28] ), .IN4(\FIFO[87][28] ), .S0(n5864), .S1(n5958), .Q(
        n5567) );
  MUX41X1 U6546 ( .IN1(\FIFO[80][28] ), .IN3(\FIFO[82][28] ), .IN2(
        \FIFO[81][28] ), .IN4(\FIFO[83][28] ), .S0(n5864), .S1(n5958), .Q(
        n5568) );
  MUX41X1 U6547 ( .IN1(n5568), .IN3(n5566), .IN2(n5567), .IN4(n5565), .S0(
        n5753), .S1(n5772), .Q(n5569) );
  MUX41X1 U6548 ( .IN1(\FIFO[76][28] ), .IN3(\FIFO[78][28] ), .IN2(
        \FIFO[77][28] ), .IN4(\FIFO[79][28] ), .S0(n5864), .S1(n5958), .Q(
        n5570) );
  MUX41X1 U6549 ( .IN1(\FIFO[72][28] ), .IN3(\FIFO[74][28] ), .IN2(
        \FIFO[73][28] ), .IN4(\FIFO[75][28] ), .S0(n5864), .S1(n5958), .Q(
        n5571) );
  MUX41X1 U6550 ( .IN1(\FIFO[68][28] ), .IN3(\FIFO[70][28] ), .IN2(
        \FIFO[69][28] ), .IN4(\FIFO[71][28] ), .S0(n5864), .S1(n5958), .Q(
        n5572) );
  MUX41X1 U6551 ( .IN1(\FIFO[64][28] ), .IN3(\FIFO[66][28] ), .IN2(
        \FIFO[65][28] ), .IN4(\FIFO[67][28] ), .S0(n5864), .S1(n5958), .Q(
        n5573) );
  MUX41X1 U6552 ( .IN1(n5573), .IN3(n5571), .IN2(n5572), .IN4(n5570), .S0(
        n5753), .S1(n5772), .Q(n5574) );
  MUX41X1 U6553 ( .IN1(n5574), .IN3(n5564), .IN2(n5569), .IN4(n5559), .S0(
        n5725), .S1(n5734), .Q(n5575) );
  MUX41X1 U6554 ( .IN1(\FIFO[60][28] ), .IN3(\FIFO[62][28] ), .IN2(
        \FIFO[61][28] ), .IN4(\FIFO[63][28] ), .S0(n5864), .S1(n5958), .Q(
        n5576) );
  MUX41X1 U6555 ( .IN1(\FIFO[56][28] ), .IN3(\FIFO[58][28] ), .IN2(
        \FIFO[57][28] ), .IN4(\FIFO[59][28] ), .S0(n5864), .S1(n5958), .Q(
        n5577) );
  MUX41X1 U6556 ( .IN1(\FIFO[52][28] ), .IN3(\FIFO[54][28] ), .IN2(
        \FIFO[53][28] ), .IN4(\FIFO[55][28] ), .S0(n5864), .S1(n5958), .Q(
        n5578) );
  MUX41X1 U6557 ( .IN1(\FIFO[48][28] ), .IN3(\FIFO[50][28] ), .IN2(
        \FIFO[49][28] ), .IN4(\FIFO[51][28] ), .S0(n5864), .S1(n5958), .Q(
        n5579) );
  MUX41X1 U6558 ( .IN1(n5579), .IN3(n5577), .IN2(n5578), .IN4(n5576), .S0(
        n5753), .S1(n5772), .Q(n5580) );
  MUX41X1 U6559 ( .IN1(\FIFO[44][28] ), .IN3(\FIFO[46][28] ), .IN2(
        \FIFO[45][28] ), .IN4(\FIFO[47][28] ), .S0(n5865), .S1(n5970), .Q(
        n5581) );
  MUX41X1 U6560 ( .IN1(\FIFO[40][28] ), .IN3(\FIFO[42][28] ), .IN2(
        \FIFO[41][28] ), .IN4(\FIFO[43][28] ), .S0(n5865), .S1(n5969), .Q(
        n5582) );
  MUX41X1 U6561 ( .IN1(\FIFO[36][28] ), .IN3(\FIFO[38][28] ), .IN2(
        \FIFO[37][28] ), .IN4(\FIFO[39][28] ), .S0(n5865), .S1(n5972), .Q(
        n5583) );
  MUX41X1 U6562 ( .IN1(\FIFO[32][28] ), .IN3(\FIFO[34][28] ), .IN2(
        \FIFO[33][28] ), .IN4(\FIFO[35][28] ), .S0(n5865), .S1(n5966), .Q(
        n5584) );
  MUX41X1 U6563 ( .IN1(n5584), .IN3(n5582), .IN2(n5583), .IN4(n5581), .S0(
        n5753), .S1(n5772), .Q(n5585) );
  MUX41X1 U6564 ( .IN1(\FIFO[28][28] ), .IN3(\FIFO[30][28] ), .IN2(
        \FIFO[29][28] ), .IN4(\FIFO[31][28] ), .S0(n5865), .S1(n5966), .Q(
        n5586) );
  MUX41X1 U6565 ( .IN1(\FIFO[24][28] ), .IN3(\FIFO[26][28] ), .IN2(
        \FIFO[25][28] ), .IN4(\FIFO[27][28] ), .S0(n5865), .S1(n5965), .Q(
        n5587) );
  MUX41X1 U6566 ( .IN1(\FIFO[20][28] ), .IN3(\FIFO[22][28] ), .IN2(
        \FIFO[21][28] ), .IN4(\FIFO[23][28] ), .S0(n5865), .S1(n5971), .Q(
        n5588) );
  MUX41X1 U6567 ( .IN1(\FIFO[16][28] ), .IN3(\FIFO[18][28] ), .IN2(
        \FIFO[17][28] ), .IN4(\FIFO[19][28] ), .S0(n5865), .S1(n5972), .Q(
        n5589) );
  MUX41X1 U6568 ( .IN1(n5589), .IN3(n5587), .IN2(n5588), .IN4(n5586), .S0(
        n5753), .S1(n5772), .Q(n5590) );
  MUX41X1 U6569 ( .IN1(\FIFO[12][28] ), .IN3(\FIFO[14][28] ), .IN2(
        \FIFO[13][28] ), .IN4(\FIFO[15][28] ), .S0(n5865), .S1(n5969), .Q(
        n5591) );
  MUX41X1 U6570 ( .IN1(\FIFO[8][28] ), .IN3(\FIFO[10][28] ), .IN2(
        \FIFO[9][28] ), .IN4(\FIFO[11][28] ), .S0(n5865), .S1(n5967), .Q(n5592) );
  MUX41X1 U6571 ( .IN1(\FIFO[4][28] ), .IN3(\FIFO[6][28] ), .IN2(\FIFO[5][28] ), .IN4(\FIFO[7][28] ), .S0(n5865), .S1(n5967), .Q(n5593) );
  MUX41X1 U6572 ( .IN1(\FIFO[0][28] ), .IN3(\FIFO[2][28] ), .IN2(\FIFO[1][28] ), .IN4(\FIFO[3][28] ), .S0(n5865), .S1(n5970), .Q(n5594) );
  MUX41X1 U6573 ( .IN1(n5594), .IN3(n5592), .IN2(n5593), .IN4(n5591), .S0(
        n5753), .S1(n5772), .Q(n5595) );
  MUX41X1 U6574 ( .IN1(n5595), .IN3(n5585), .IN2(n5590), .IN4(n5580), .S0(
        n5727), .S1(n5734), .Q(n5596) );
  MUX21X1 U6575 ( .IN1(n5596), .IN2(n5575), .S(n5724), .Q(N222) );
  MUX41X1 U6576 ( .IN1(\FIFO[124][29] ), .IN3(\FIFO[126][29] ), .IN2(
        \FIFO[125][29] ), .IN4(\FIFO[127][29] ), .S0(n5866), .S1(n5959), .Q(
        n5597) );
  MUX41X1 U6577 ( .IN1(\FIFO[120][29] ), .IN3(\FIFO[122][29] ), .IN2(
        \FIFO[121][29] ), .IN4(\FIFO[123][29] ), .S0(n5866), .S1(n5959), .Q(
        n5598) );
  MUX41X1 U6578 ( .IN1(\FIFO[116][29] ), .IN3(\FIFO[118][29] ), .IN2(
        \FIFO[117][29] ), .IN4(\FIFO[119][29] ), .S0(n5866), .S1(n5959), .Q(
        n5599) );
  MUX41X1 U6579 ( .IN1(\FIFO[112][29] ), .IN3(\FIFO[114][29] ), .IN2(
        \FIFO[113][29] ), .IN4(\FIFO[115][29] ), .S0(n5866), .S1(n5959), .Q(
        n5600) );
  MUX41X1 U6580 ( .IN1(n5600), .IN3(n5598), .IN2(n5599), .IN4(n5597), .S0(
        n5754), .S1(n5773), .Q(n5601) );
  MUX41X1 U6581 ( .IN1(\FIFO[108][29] ), .IN3(\FIFO[110][29] ), .IN2(
        \FIFO[109][29] ), .IN4(\FIFO[111][29] ), .S0(n5866), .S1(n5959), .Q(
        n5602) );
  MUX41X1 U6582 ( .IN1(\FIFO[104][29] ), .IN3(\FIFO[106][29] ), .IN2(
        \FIFO[105][29] ), .IN4(\FIFO[107][29] ), .S0(n5866), .S1(n5959), .Q(
        n5603) );
  MUX41X1 U6583 ( .IN1(\FIFO[100][29] ), .IN3(\FIFO[102][29] ), .IN2(
        \FIFO[101][29] ), .IN4(\FIFO[103][29] ), .S0(n5866), .S1(n5959), .Q(
        n5604) );
  MUX41X1 U6584 ( .IN1(\FIFO[96][29] ), .IN3(\FIFO[98][29] ), .IN2(
        \FIFO[97][29] ), .IN4(\FIFO[99][29] ), .S0(n5866), .S1(n5959), .Q(
        n5605) );
  MUX41X1 U6585 ( .IN1(n5605), .IN3(n5603), .IN2(n5604), .IN4(n5602), .S0(
        n5754), .S1(n5773), .Q(n5606) );
  MUX41X1 U6586 ( .IN1(\FIFO[92][29] ), .IN3(\FIFO[94][29] ), .IN2(
        \FIFO[93][29] ), .IN4(\FIFO[95][29] ), .S0(n5866), .S1(n5959), .Q(
        n5607) );
  MUX41X1 U6587 ( .IN1(\FIFO[88][29] ), .IN3(\FIFO[90][29] ), .IN2(
        \FIFO[89][29] ), .IN4(\FIFO[91][29] ), .S0(n5866), .S1(n5959), .Q(
        n5608) );
  MUX41X1 U6588 ( .IN1(\FIFO[84][29] ), .IN3(\FIFO[86][29] ), .IN2(
        \FIFO[85][29] ), .IN4(\FIFO[87][29] ), .S0(n5866), .S1(n5959), .Q(
        n5609) );
  MUX41X1 U6589 ( .IN1(\FIFO[80][29] ), .IN3(\FIFO[82][29] ), .IN2(
        \FIFO[81][29] ), .IN4(\FIFO[83][29] ), .S0(n5866), .S1(n5959), .Q(
        n5610) );
  MUX41X1 U6590 ( .IN1(n5610), .IN3(n5608), .IN2(n5609), .IN4(n5607), .S0(
        n5754), .S1(n5773), .Q(n5611) );
  MUX41X1 U6591 ( .IN1(\FIFO[76][29] ), .IN3(\FIFO[78][29] ), .IN2(
        \FIFO[77][29] ), .IN4(\FIFO[79][29] ), .S0(n5867), .S1(n5960), .Q(
        n5612) );
  MUX41X1 U6592 ( .IN1(\FIFO[72][29] ), .IN3(\FIFO[74][29] ), .IN2(
        \FIFO[73][29] ), .IN4(\FIFO[75][29] ), .S0(n5867), .S1(n5960), .Q(
        n5613) );
  MUX41X1 U6593 ( .IN1(\FIFO[68][29] ), .IN3(\FIFO[70][29] ), .IN2(
        \FIFO[69][29] ), .IN4(\FIFO[71][29] ), .S0(n5867), .S1(n5960), .Q(
        n5614) );
  MUX41X1 U6594 ( .IN1(\FIFO[64][29] ), .IN3(\FIFO[66][29] ), .IN2(
        \FIFO[65][29] ), .IN4(\FIFO[67][29] ), .S0(n5867), .S1(n5960), .Q(
        n5615) );
  MUX41X1 U6595 ( .IN1(n5615), .IN3(n5613), .IN2(n5614), .IN4(n5612), .S0(
        n5754), .S1(n5773), .Q(n5616) );
  MUX41X1 U6596 ( .IN1(n5616), .IN3(n5606), .IN2(n5611), .IN4(n5601), .S0(
        n5725), .S1(n5734), .Q(n5617) );
  MUX41X1 U6597 ( .IN1(\FIFO[60][29] ), .IN3(\FIFO[62][29] ), .IN2(
        \FIFO[61][29] ), .IN4(\FIFO[63][29] ), .S0(n5867), .S1(n5960), .Q(
        n5618) );
  MUX41X1 U6598 ( .IN1(\FIFO[56][29] ), .IN3(\FIFO[58][29] ), .IN2(
        \FIFO[57][29] ), .IN4(\FIFO[59][29] ), .S0(n5867), .S1(n5960), .Q(
        n5619) );
  MUX41X1 U6599 ( .IN1(\FIFO[52][29] ), .IN3(\FIFO[54][29] ), .IN2(
        \FIFO[53][29] ), .IN4(\FIFO[55][29] ), .S0(n5867), .S1(n5960), .Q(
        n5620) );
  MUX41X1 U6600 ( .IN1(\FIFO[48][29] ), .IN3(\FIFO[50][29] ), .IN2(
        \FIFO[49][29] ), .IN4(\FIFO[51][29] ), .S0(n5867), .S1(n5960), .Q(
        n5621) );
  MUX41X1 U6601 ( .IN1(n5621), .IN3(n5619), .IN2(n5620), .IN4(n5618), .S0(
        n5754), .S1(n5773), .Q(n5622) );
  MUX41X1 U6602 ( .IN1(\FIFO[44][29] ), .IN3(\FIFO[46][29] ), .IN2(
        \FIFO[45][29] ), .IN4(\FIFO[47][29] ), .S0(n5867), .S1(n5960), .Q(
        n5623) );
  MUX41X1 U6603 ( .IN1(\FIFO[40][29] ), .IN3(\FIFO[42][29] ), .IN2(
        \FIFO[41][29] ), .IN4(\FIFO[43][29] ), .S0(n5867), .S1(n5960), .Q(
        n5624) );
  MUX41X1 U6604 ( .IN1(\FIFO[36][29] ), .IN3(\FIFO[38][29] ), .IN2(
        \FIFO[37][29] ), .IN4(\FIFO[39][29] ), .S0(n5867), .S1(n5960), .Q(
        n5625) );
  MUX41X1 U6605 ( .IN1(\FIFO[32][29] ), .IN3(\FIFO[34][29] ), .IN2(
        \FIFO[33][29] ), .IN4(\FIFO[35][29] ), .S0(n5867), .S1(n5960), .Q(
        n5626) );
  MUX41X1 U6606 ( .IN1(n5626), .IN3(n5624), .IN2(n5625), .IN4(n5623), .S0(
        n5754), .S1(n5773), .Q(n5627) );
  MUX41X1 U6607 ( .IN1(\FIFO[28][29] ), .IN3(\FIFO[30][29] ), .IN2(
        \FIFO[29][29] ), .IN4(\FIFO[31][29] ), .S0(n5868), .S1(n5961), .Q(
        n5628) );
  MUX41X1 U6608 ( .IN1(\FIFO[24][29] ), .IN3(\FIFO[26][29] ), .IN2(
        \FIFO[25][29] ), .IN4(\FIFO[27][29] ), .S0(n5868), .S1(n5961), .Q(
        n5629) );
  MUX41X1 U6609 ( .IN1(\FIFO[20][29] ), .IN3(\FIFO[22][29] ), .IN2(
        \FIFO[21][29] ), .IN4(\FIFO[23][29] ), .S0(n5868), .S1(n5961), .Q(
        n5630) );
  MUX41X1 U6610 ( .IN1(\FIFO[16][29] ), .IN3(\FIFO[18][29] ), .IN2(
        \FIFO[17][29] ), .IN4(\FIFO[19][29] ), .S0(n5868), .S1(n5961), .Q(
        n5631) );
  MUX41X1 U6611 ( .IN1(n5631), .IN3(n5629), .IN2(n5630), .IN4(n5628), .S0(
        n5754), .S1(n5773), .Q(n5632) );
  MUX41X1 U6612 ( .IN1(\FIFO[12][29] ), .IN3(\FIFO[14][29] ), .IN2(
        \FIFO[13][29] ), .IN4(\FIFO[15][29] ), .S0(n5868), .S1(n5961), .Q(
        n5633) );
  MUX41X1 U6613 ( .IN1(\FIFO[8][29] ), .IN3(\FIFO[10][29] ), .IN2(
        \FIFO[9][29] ), .IN4(\FIFO[11][29] ), .S0(n5868), .S1(n5961), .Q(n5634) );
  MUX41X1 U6614 ( .IN1(\FIFO[4][29] ), .IN3(\FIFO[6][29] ), .IN2(\FIFO[5][29] ), .IN4(\FIFO[7][29] ), .S0(n5868), .S1(n5961), .Q(n5635) );
  MUX41X1 U6615 ( .IN1(\FIFO[0][29] ), .IN3(\FIFO[2][29] ), .IN2(\FIFO[1][29] ), .IN4(\FIFO[3][29] ), .S0(n5868), .S1(n5961), .Q(n5636) );
  MUX41X1 U6616 ( .IN1(n5636), .IN3(n5634), .IN2(n5635), .IN4(n5633), .S0(
        n5754), .S1(n5773), .Q(n5637) );
  MUX41X1 U6617 ( .IN1(n5637), .IN3(n5627), .IN2(n5632), .IN4(n5622), .S0(
        n5728), .S1(n5734), .Q(n5638) );
  MUX21X1 U6618 ( .IN1(n5638), .IN2(n5617), .S(n5724), .Q(N221) );
  MUX41X1 U6619 ( .IN1(\FIFO[124][30] ), .IN3(\FIFO[126][30] ), .IN2(
        \FIFO[125][30] ), .IN4(\FIFO[127][30] ), .S0(n5868), .S1(n5961), .Q(
        n5639) );
  MUX41X1 U6620 ( .IN1(\FIFO[120][30] ), .IN3(\FIFO[122][30] ), .IN2(
        \FIFO[121][30] ), .IN4(\FIFO[123][30] ), .S0(n5868), .S1(n5961), .Q(
        n5640) );
  MUX41X1 U6621 ( .IN1(\FIFO[116][30] ), .IN3(\FIFO[118][30] ), .IN2(
        \FIFO[117][30] ), .IN4(\FIFO[119][30] ), .S0(n5868), .S1(n5961), .Q(
        n5641) );
  MUX41X1 U6622 ( .IN1(\FIFO[112][30] ), .IN3(\FIFO[114][30] ), .IN2(
        \FIFO[113][30] ), .IN4(\FIFO[115][30] ), .S0(n5868), .S1(n5961), .Q(
        n5642) );
  MUX41X1 U6623 ( .IN1(n5642), .IN3(n5640), .IN2(n5641), .IN4(n5639), .S0(
        n5754), .S1(n5773), .Q(n5643) );
  MUX41X1 U6624 ( .IN1(\FIFO[108][30] ), .IN3(\FIFO[110][30] ), .IN2(
        \FIFO[109][30] ), .IN4(\FIFO[111][30] ), .S0(n5869), .S1(n5962), .Q(
        n5644) );
  MUX41X1 U6625 ( .IN1(\FIFO[104][30] ), .IN3(\FIFO[106][30] ), .IN2(
        \FIFO[105][30] ), .IN4(\FIFO[107][30] ), .S0(n5869), .S1(n5962), .Q(
        n5645) );
  MUX41X1 U6626 ( .IN1(\FIFO[100][30] ), .IN3(\FIFO[102][30] ), .IN2(
        \FIFO[101][30] ), .IN4(\FIFO[103][30] ), .S0(n5869), .S1(n5962), .Q(
        n5646) );
  MUX41X1 U6627 ( .IN1(\FIFO[96][30] ), .IN3(\FIFO[98][30] ), .IN2(
        \FIFO[97][30] ), .IN4(\FIFO[99][30] ), .S0(n5869), .S1(n5962), .Q(
        n5647) );
  MUX41X1 U6628 ( .IN1(n5647), .IN3(n5645), .IN2(n5646), .IN4(n5644), .S0(
        n5754), .S1(n5773), .Q(n5648) );
  MUX41X1 U6629 ( .IN1(\FIFO[92][30] ), .IN3(\FIFO[94][30] ), .IN2(
        \FIFO[93][30] ), .IN4(\FIFO[95][30] ), .S0(n5869), .S1(n5962), .Q(
        n5649) );
  MUX41X1 U6630 ( .IN1(\FIFO[88][30] ), .IN3(\FIFO[90][30] ), .IN2(
        \FIFO[89][30] ), .IN4(\FIFO[91][30] ), .S0(n5869), .S1(n5962), .Q(
        n5650) );
  MUX41X1 U6631 ( .IN1(\FIFO[84][30] ), .IN3(\FIFO[86][30] ), .IN2(
        \FIFO[85][30] ), .IN4(\FIFO[87][30] ), .S0(n5869), .S1(n5962), .Q(
        n5651) );
  MUX41X1 U6632 ( .IN1(\FIFO[80][30] ), .IN3(\FIFO[82][30] ), .IN2(
        \FIFO[81][30] ), .IN4(\FIFO[83][30] ), .S0(n5869), .S1(n5962), .Q(
        n5652) );
  MUX41X1 U6633 ( .IN1(n5652), .IN3(n5650), .IN2(n5651), .IN4(n5649), .S0(
        n5754), .S1(n5773), .Q(n5653) );
  MUX41X1 U6634 ( .IN1(\FIFO[76][30] ), .IN3(\FIFO[78][30] ), .IN2(
        \FIFO[77][30] ), .IN4(\FIFO[79][30] ), .S0(n5869), .S1(n5962), .Q(
        n5654) );
  MUX41X1 U6635 ( .IN1(\FIFO[72][30] ), .IN3(\FIFO[74][30] ), .IN2(
        \FIFO[73][30] ), .IN4(\FIFO[75][30] ), .S0(n5869), .S1(n5962), .Q(
        n5655) );
  MUX41X1 U6636 ( .IN1(\FIFO[68][30] ), .IN3(\FIFO[70][30] ), .IN2(
        \FIFO[69][30] ), .IN4(\FIFO[71][30] ), .S0(n5869), .S1(n5962), .Q(
        n5656) );
  MUX41X1 U6637 ( .IN1(\FIFO[64][30] ), .IN3(\FIFO[66][30] ), .IN2(
        \FIFO[65][30] ), .IN4(\FIFO[67][30] ), .S0(n5869), .S1(n5962), .Q(
        n5657) );
  MUX41X1 U6638 ( .IN1(n5657), .IN3(n5655), .IN2(n5656), .IN4(n5654), .S0(
        n5754), .S1(n5773), .Q(n5658) );
  MUX41X1 U6639 ( .IN1(n5658), .IN3(n5648), .IN2(n5653), .IN4(n5643), .S0(
        n5725), .S1(n5734), .Q(n5659) );
  MUX41X1 U6640 ( .IN1(\FIFO[60][30] ), .IN3(\FIFO[62][30] ), .IN2(
        \FIFO[61][30] ), .IN4(\FIFO[63][30] ), .S0(n5870), .S1(n5963), .Q(
        n5660) );
  MUX41X1 U6641 ( .IN1(\FIFO[56][30] ), .IN3(\FIFO[58][30] ), .IN2(
        \FIFO[57][30] ), .IN4(\FIFO[59][30] ), .S0(n5870), .S1(n5963), .Q(
        n5661) );
  MUX41X1 U6642 ( .IN1(\FIFO[52][30] ), .IN3(\FIFO[54][30] ), .IN2(
        \FIFO[53][30] ), .IN4(\FIFO[55][30] ), .S0(n5870), .S1(n5963), .Q(
        n5662) );
  MUX41X1 U6643 ( .IN1(\FIFO[48][30] ), .IN3(\FIFO[50][30] ), .IN2(
        \FIFO[49][30] ), .IN4(\FIFO[51][30] ), .S0(n5870), .S1(n5963), .Q(
        n5663) );
  MUX41X1 U6644 ( .IN1(n5663), .IN3(n5661), .IN2(n5662), .IN4(n5660), .S0(
        n5755), .S1(n5774), .Q(n5664) );
  MUX41X1 U6645 ( .IN1(\FIFO[44][30] ), .IN3(\FIFO[46][30] ), .IN2(
        \FIFO[45][30] ), .IN4(\FIFO[47][30] ), .S0(n5870), .S1(n5963), .Q(
        n5665) );
  MUX41X1 U6646 ( .IN1(\FIFO[40][30] ), .IN3(\FIFO[42][30] ), .IN2(
        \FIFO[41][30] ), .IN4(\FIFO[43][30] ), .S0(n5870), .S1(n5963), .Q(
        n5666) );
  MUX41X1 U6647 ( .IN1(\FIFO[36][30] ), .IN3(\FIFO[38][30] ), .IN2(
        \FIFO[37][30] ), .IN4(\FIFO[39][30] ), .S0(n5870), .S1(n5963), .Q(
        n5667) );
  MUX41X1 U6648 ( .IN1(\FIFO[32][30] ), .IN3(\FIFO[34][30] ), .IN2(
        \FIFO[33][30] ), .IN4(\FIFO[35][30] ), .S0(n5870), .S1(n5963), .Q(
        n5668) );
  MUX41X1 U6649 ( .IN1(n5668), .IN3(n5666), .IN2(n5667), .IN4(n5665), .S0(
        n5755), .S1(n5774), .Q(n5669) );
  MUX41X1 U6650 ( .IN1(\FIFO[28][30] ), .IN3(\FIFO[30][30] ), .IN2(
        \FIFO[29][30] ), .IN4(\FIFO[31][30] ), .S0(n5870), .S1(n5963), .Q(
        n5670) );
  MUX41X1 U6651 ( .IN1(\FIFO[24][30] ), .IN3(\FIFO[26][30] ), .IN2(
        \FIFO[25][30] ), .IN4(\FIFO[27][30] ), .S0(n5870), .S1(n5963), .Q(
        n5671) );
  MUX41X1 U6652 ( .IN1(\FIFO[20][30] ), .IN3(\FIFO[22][30] ), .IN2(
        \FIFO[21][30] ), .IN4(\FIFO[23][30] ), .S0(n5870), .S1(n5963), .Q(
        n5672) );
  MUX41X1 U6653 ( .IN1(\FIFO[16][30] ), .IN3(\FIFO[18][30] ), .IN2(
        \FIFO[17][30] ), .IN4(\FIFO[19][30] ), .S0(n5870), .S1(n5963), .Q(
        n5673) );
  MUX41X1 U6654 ( .IN1(n5673), .IN3(n5671), .IN2(n5672), .IN4(n5670), .S0(
        n5755), .S1(n5774), .Q(n5674) );
  MUX41X1 U6655 ( .IN1(\FIFO[12][30] ), .IN3(\FIFO[14][30] ), .IN2(
        \FIFO[13][30] ), .IN4(\FIFO[15][30] ), .S0(n5871), .S1(n5964), .Q(
        n5675) );
  MUX41X1 U6656 ( .IN1(\FIFO[8][30] ), .IN3(\FIFO[10][30] ), .IN2(
        \FIFO[9][30] ), .IN4(\FIFO[11][30] ), .S0(n5871), .S1(n5964), .Q(n5676) );
  MUX41X1 U6657 ( .IN1(\FIFO[4][30] ), .IN3(\FIFO[6][30] ), .IN2(\FIFO[5][30] ), .IN4(\FIFO[7][30] ), .S0(n5871), .S1(n5964), .Q(n5677) );
  MUX41X1 U6658 ( .IN1(\FIFO[0][30] ), .IN3(\FIFO[2][30] ), .IN2(\FIFO[1][30] ), .IN4(\FIFO[3][30] ), .S0(n5871), .S1(n5964), .Q(n5678) );
  MUX41X1 U6659 ( .IN1(n5678), .IN3(n5676), .IN2(n5677), .IN4(n5675), .S0(
        n5755), .S1(n5774), .Q(n5679) );
  MUX41X1 U6660 ( .IN1(n5679), .IN3(n5669), .IN2(n5674), .IN4(n5664), .S0(
        n5725), .S1(n5734), .Q(n5680) );
  MUX21X1 U6661 ( .IN1(n5680), .IN2(n5659), .S(n5724), .Q(N220) );
  MUX41X1 U6662 ( .IN1(\FIFO[124][31] ), .IN3(\FIFO[126][31] ), .IN2(
        \FIFO[125][31] ), .IN4(\FIFO[127][31] ), .S0(n5871), .S1(n5964), .Q(
        n5681) );
  MUX41X1 U6663 ( .IN1(\FIFO[120][31] ), .IN3(\FIFO[122][31] ), .IN2(
        \FIFO[121][31] ), .IN4(\FIFO[123][31] ), .S0(n5871), .S1(n5964), .Q(
        n5682) );
  MUX41X1 U6664 ( .IN1(\FIFO[116][31] ), .IN3(\FIFO[118][31] ), .IN2(
        \FIFO[117][31] ), .IN4(\FIFO[119][31] ), .S0(n5871), .S1(n5964), .Q(
        n5683) );
  MUX41X1 U6665 ( .IN1(\FIFO[112][31] ), .IN3(\FIFO[114][31] ), .IN2(
        \FIFO[113][31] ), .IN4(\FIFO[115][31] ), .S0(n5871), .S1(n5964), .Q(
        n5684) );
  MUX41X1 U6666 ( .IN1(n5684), .IN3(n5682), .IN2(n5683), .IN4(n5681), .S0(
        n5755), .S1(n5774), .Q(n5685) );
  MUX41X1 U6667 ( .IN1(\FIFO[108][31] ), .IN3(\FIFO[110][31] ), .IN2(
        \FIFO[109][31] ), .IN4(\FIFO[111][31] ), .S0(n5871), .S1(n5964), .Q(
        n5686) );
  MUX41X1 U6668 ( .IN1(\FIFO[104][31] ), .IN3(\FIFO[106][31] ), .IN2(
        \FIFO[105][31] ), .IN4(\FIFO[107][31] ), .S0(n5871), .S1(n5964), .Q(
        n5687) );
  MUX41X1 U6669 ( .IN1(\FIFO[100][31] ), .IN3(\FIFO[102][31] ), .IN2(
        \FIFO[101][31] ), .IN4(\FIFO[103][31] ), .S0(n5871), .S1(n5964), .Q(
        n5688) );
  MUX41X1 U6670 ( .IN1(\FIFO[96][31] ), .IN3(\FIFO[98][31] ), .IN2(
        \FIFO[97][31] ), .IN4(\FIFO[99][31] ), .S0(n5871), .S1(n5964), .Q(
        n5689) );
  MUX41X1 U6671 ( .IN1(n5689), .IN3(n5687), .IN2(n5688), .IN4(n5686), .S0(
        n5755), .S1(n5774), .Q(n5690) );
  MUX41X1 U6672 ( .IN1(\FIFO[92][31] ), .IN3(\FIFO[94][31] ), .IN2(
        \FIFO[93][31] ), .IN4(\FIFO[95][31] ), .S0(n5872), .S1(n5895), .Q(
        n5691) );
  MUX41X1 U6673 ( .IN1(\FIFO[88][31] ), .IN3(\FIFO[90][31] ), .IN2(
        \FIFO[89][31] ), .IN4(\FIFO[91][31] ), .S0(n5872), .S1(n5890), .Q(
        n5692) );
  MUX41X1 U6674 ( .IN1(\FIFO[84][31] ), .IN3(\FIFO[86][31] ), .IN2(
        \FIFO[85][31] ), .IN4(\FIFO[87][31] ), .S0(n5872), .S1(n5877), .Q(
        n5693) );
  MUX41X1 U6675 ( .IN1(\FIFO[80][31] ), .IN3(\FIFO[82][31] ), .IN2(
        \FIFO[81][31] ), .IN4(\FIFO[83][31] ), .S0(n5872), .S1(n5875), .Q(
        n5694) );
  MUX41X1 U6676 ( .IN1(n5694), .IN3(n5692), .IN2(n5693), .IN4(n5691), .S0(
        n5755), .S1(n5774), .Q(n5695) );
  MUX41X1 U6677 ( .IN1(\FIFO[76][31] ), .IN3(\FIFO[78][31] ), .IN2(
        \FIFO[77][31] ), .IN4(\FIFO[79][31] ), .S0(n5872), .S1(n5891), .Q(
        n5696) );
  MUX41X1 U6678 ( .IN1(\FIFO[72][31] ), .IN3(\FIFO[74][31] ), .IN2(
        \FIFO[73][31] ), .IN4(\FIFO[75][31] ), .S0(n5872), .S1(n5971), .Q(
        n5697) );
  MUX41X1 U6679 ( .IN1(\FIFO[68][31] ), .IN3(\FIFO[70][31] ), .IN2(
        \FIFO[69][31] ), .IN4(\FIFO[71][31] ), .S0(n5872), .S1(n5880), .Q(
        n5698) );
  MUX41X1 U6680 ( .IN1(\FIFO[64][31] ), .IN3(\FIFO[66][31] ), .IN2(
        \FIFO[65][31] ), .IN4(\FIFO[67][31] ), .S0(n5872), .S1(n5879), .Q(
        n5699) );
  MUX41X1 U6681 ( .IN1(n5699), .IN3(n5697), .IN2(n5698), .IN4(n5696), .S0(
        n5755), .S1(n5774), .Q(n5700) );
  MUX41X1 U6682 ( .IN1(n5700), .IN3(n5690), .IN2(n5695), .IN4(n5685), .S0(
        n5725), .S1(n5734), .Q(n5701) );
  MUX41X1 U6683 ( .IN1(\FIFO[60][31] ), .IN3(\FIFO[62][31] ), .IN2(
        \FIFO[61][31] ), .IN4(\FIFO[63][31] ), .S0(n5872), .S1(n5876), .Q(
        n5702) );
  MUX41X1 U6684 ( .IN1(\FIFO[56][31] ), .IN3(\FIFO[58][31] ), .IN2(
        \FIFO[57][31] ), .IN4(\FIFO[59][31] ), .S0(n5872), .S1(n5882), .Q(
        n5703) );
  MUX41X1 U6685 ( .IN1(\FIFO[52][31] ), .IN3(\FIFO[54][31] ), .IN2(
        \FIFO[53][31] ), .IN4(\FIFO[55][31] ), .S0(n5872), .S1(n5965), .Q(
        n5704) );
  MUX41X1 U6686 ( .IN1(\FIFO[48][31] ), .IN3(\FIFO[50][31] ), .IN2(
        \FIFO[49][31] ), .IN4(\FIFO[51][31] ), .S0(n5872), .S1(n5874), .Q(
        n5705) );
  MUX41X1 U6687 ( .IN1(n5705), .IN3(n5703), .IN2(n5704), .IN4(n5702), .S0(
        n5755), .S1(n5774), .Q(n5706) );
  MUX41X1 U6688 ( .IN1(\FIFO[44][31] ), .IN3(\FIFO[46][31] ), .IN2(
        \FIFO[45][31] ), .IN4(\FIFO[47][31] ), .S0(n5873), .S1(n5970), .Q(
        n5707) );
  MUX41X1 U6689 ( .IN1(\FIFO[40][31] ), .IN3(\FIFO[42][31] ), .IN2(
        \FIFO[41][31] ), .IN4(\FIFO[43][31] ), .S0(n5873), .S1(n5969), .Q(
        n5708) );
  MUX41X1 U6690 ( .IN1(\FIFO[36][31] ), .IN3(\FIFO[38][31] ), .IN2(
        \FIFO[37][31] ), .IN4(\FIFO[39][31] ), .S0(n5873), .S1(n5876), .Q(
        n5709) );
  MUX41X1 U6691 ( .IN1(\FIFO[32][31] ), .IN3(\FIFO[34][31] ), .IN2(
        \FIFO[33][31] ), .IN4(\FIFO[35][31] ), .S0(n5873), .S1(n5875), .Q(
        n5710) );
  MUX41X1 U6692 ( .IN1(n5710), .IN3(n5708), .IN2(n5709), .IN4(n5707), .S0(
        n5755), .S1(n5774), .Q(n5711) );
  MUX41X1 U6693 ( .IN1(\FIFO[28][31] ), .IN3(\FIFO[30][31] ), .IN2(
        \FIFO[29][31] ), .IN4(\FIFO[31][31] ), .S0(n5873), .S1(n5966), .Q(
        n5712) );
  MUX41X1 U6694 ( .IN1(\FIFO[24][31] ), .IN3(\FIFO[26][31] ), .IN2(
        \FIFO[25][31] ), .IN4(\FIFO[27][31] ), .S0(n5873), .S1(n5877), .Q(
        n5713) );
  MUX41X1 U6695 ( .IN1(\FIFO[20][31] ), .IN3(\FIFO[22][31] ), .IN2(
        \FIFO[21][31] ), .IN4(\FIFO[23][31] ), .S0(n5873), .S1(n5970), .Q(
        n5714) );
  MUX41X1 U6696 ( .IN1(\FIFO[16][31] ), .IN3(\FIFO[18][31] ), .IN2(
        \FIFO[17][31] ), .IN4(\FIFO[19][31] ), .S0(n5873), .S1(n5969), .Q(
        n5715) );
  MUX41X1 U6697 ( .IN1(n5715), .IN3(n5713), .IN2(n5714), .IN4(n5712), .S0(
        n5755), .S1(n5774), .Q(n5716) );
  MUX41X1 U6698 ( .IN1(\FIFO[12][31] ), .IN3(\FIFO[14][31] ), .IN2(
        \FIFO[13][31] ), .IN4(\FIFO[15][31] ), .S0(n5873), .S1(n5968), .Q(
        n5717) );
  MUX41X1 U6699 ( .IN1(\FIFO[8][31] ), .IN3(\FIFO[10][31] ), .IN2(
        \FIFO[9][31] ), .IN4(\FIFO[11][31] ), .S0(n5873), .S1(n5971), .Q(n5718) );
  MUX41X1 U6700 ( .IN1(\FIFO[4][31] ), .IN3(\FIFO[6][31] ), .IN2(\FIFO[5][31] ), .IN4(\FIFO[7][31] ), .S0(n5873), .S1(n5972), .Q(n5719) );
  MUX41X1 U6701 ( .IN1(\FIFO[0][31] ), .IN3(\FIFO[2][31] ), .IN2(\FIFO[1][31] ), .IN4(\FIFO[3][31] ), .S0(n5873), .S1(n5967), .Q(n5720) );
  MUX41X1 U6702 ( .IN1(n5720), .IN3(n5718), .IN2(n5719), .IN4(n5717), .S0(
        n5755), .S1(n5774), .Q(n5721) );
  MUX41X1 U6703 ( .IN1(n5721), .IN3(n5711), .IN2(n5716), .IN4(n5706), .S0(
        n5729), .S1(n5734), .Q(n5722) );
  MUX21X1 U6704 ( .IN1(n5722), .IN2(n5701), .S(n5724), .Q(N219) );
  NBUFFX4 U6705 ( .INP(n5779), .Z(n5759) );
  NBUFFX4 U6706 ( .INP(n5777), .Z(n5760) );
  NBUFFX4 U6707 ( .INP(n5777), .Z(n5761) );
  NBUFFX4 U6708 ( .INP(n5777), .Z(n5762) );
  NBUFFX4 U6709 ( .INP(n5778), .Z(n5763) );
  NBUFFX4 U6710 ( .INP(n5778), .Z(n5764) );
  NBUFFX4 U6711 ( .INP(n5778), .Z(n5765) );
  NBUFFX4 U6712 ( .INP(n5779), .Z(n5766) );
  NBUFFX4 U6713 ( .INP(n5779), .Z(n5767) );
  NBUFFX4 U6714 ( .INP(n5779), .Z(n5768) );
  NBUFFX4 U6715 ( .INP(n5780), .Z(n5769) );
  NBUFFX4 U6716 ( .INP(n5780), .Z(n5770) );
  NBUFFX4 U6717 ( .INP(n5780), .Z(n5771) );
  NBUFFX4 U6718 ( .INP(n5781), .Z(n5772) );
  NBUFFX4 U6719 ( .INP(n5781), .Z(n5773) );
  NBUFFX4 U6720 ( .INP(n5781), .Z(n5774) );
  NBUFFX4 U6721 ( .INP(n5896), .Z(n5897) );
  NBUFFX4 U6722 ( .INP(n5896), .Z(n5898) );
  NBUFFX4 U6723 ( .INP(n5896), .Z(n5899) );
  NBUFFX4 U6724 ( .INP(n5895), .Z(n5900) );
  NBUFFX4 U6725 ( .INP(n5895), .Z(n5901) );
  NBUFFX4 U6726 ( .INP(n5895), .Z(n5902) );
  NBUFFX4 U6727 ( .INP(n5894), .Z(n5903) );
  NBUFFX4 U6728 ( .INP(n5894), .Z(n5904) );
  NBUFFX4 U6729 ( .INP(n5894), .Z(n5905) );
  NBUFFX4 U6730 ( .INP(n5893), .Z(n5906) );
  NBUFFX4 U6731 ( .INP(n5893), .Z(n5907) );
  NBUFFX4 U6732 ( .INP(n5893), .Z(n5908) );
  NBUFFX4 U6733 ( .INP(n5892), .Z(n5909) );
  NBUFFX4 U6734 ( .INP(n5892), .Z(n5910) );
  NBUFFX4 U6735 ( .INP(n5892), .Z(n5911) );
  NBUFFX4 U6736 ( .INP(n5891), .Z(n5912) );
  NBUFFX4 U6737 ( .INP(n5891), .Z(n5913) );
  NBUFFX4 U6738 ( .INP(n5891), .Z(n5914) );
  NBUFFX4 U6739 ( .INP(n5890), .Z(n5915) );
  NBUFFX4 U6740 ( .INP(n5890), .Z(n5916) );
  NBUFFX4 U6741 ( .INP(n5890), .Z(n5917) );
  NBUFFX4 U6742 ( .INP(n5889), .Z(n5918) );
  NBUFFX4 U6743 ( .INP(n5889), .Z(n5919) );
  NBUFFX4 U6744 ( .INP(n5889), .Z(n5920) );
  NBUFFX4 U6745 ( .INP(n5888), .Z(n5921) );
  NBUFFX4 U6746 ( .INP(n5888), .Z(n5922) );
  NBUFFX4 U6747 ( .INP(n5888), .Z(n5923) );
  NBUFFX4 U6748 ( .INP(n5887), .Z(n5924) );
  NBUFFX4 U6749 ( .INP(n5887), .Z(n5925) );
  NBUFFX4 U6750 ( .INP(n5887), .Z(n5926) );
  NBUFFX4 U6751 ( .INP(n5886), .Z(n5927) );
  NBUFFX4 U6752 ( .INP(n5886), .Z(n5928) );
  NBUFFX4 U6753 ( .INP(n5886), .Z(n5929) );
  NBUFFX4 U6754 ( .INP(n5885), .Z(n5930) );
  NBUFFX4 U6755 ( .INP(n5885), .Z(n5931) );
  NBUFFX4 U6756 ( .INP(n5885), .Z(n5932) );
  NBUFFX4 U6757 ( .INP(n5884), .Z(n5933) );
  NBUFFX4 U6758 ( .INP(n5884), .Z(n5934) );
  NBUFFX4 U6759 ( .INP(n5884), .Z(n5935) );
  NBUFFX4 U6760 ( .INP(n5883), .Z(n5936) );
  NBUFFX4 U6761 ( .INP(n5883), .Z(n5937) );
  NBUFFX4 U6762 ( .INP(n5883), .Z(n5938) );
  NBUFFX4 U6763 ( .INP(n5882), .Z(n5939) );
  NBUFFX4 U6764 ( .INP(n5882), .Z(n5940) );
  NBUFFX4 U6765 ( .INP(n5882), .Z(n5941) );
  NBUFFX4 U6766 ( .INP(n5881), .Z(n5942) );
  NBUFFX4 U6767 ( .INP(n5881), .Z(n5943) );
  NBUFFX4 U6768 ( .INP(n5881), .Z(n5944) );
  NBUFFX4 U6769 ( .INP(n5880), .Z(n5945) );
  NBUFFX4 U6770 ( .INP(n5880), .Z(n5946) );
  NBUFFX4 U6771 ( .INP(n5880), .Z(n5947) );
  NBUFFX4 U6772 ( .INP(n5879), .Z(n5948) );
  NBUFFX4 U6773 ( .INP(n5879), .Z(n5949) );
  NBUFFX4 U6774 ( .INP(n5879), .Z(n5950) );
  NBUFFX4 U6775 ( .INP(n5878), .Z(n5951) );
  NBUFFX4 U6776 ( .INP(n5878), .Z(n5952) );
  NBUFFX4 U6777 ( .INP(n5878), .Z(n5953) );
  NBUFFX4 U6778 ( .INP(n5877), .Z(n5954) );
  NBUFFX4 U6779 ( .INP(n5877), .Z(n5955) );
  NBUFFX4 U6780 ( .INP(n5877), .Z(n5956) );
  NBUFFX4 U6781 ( .INP(n5876), .Z(n5957) );
  NBUFFX4 U6782 ( .INP(n5876), .Z(n5958) );
  NBUFFX4 U6783 ( .INP(n5875), .Z(n5959) );
  NBUFFX4 U6784 ( .INP(n5875), .Z(n5960) );
  NBUFFX4 U6785 ( .INP(n5875), .Z(n5961) );
  NBUFFX4 U6786 ( .INP(n5874), .Z(n5962) );
  NBUFFX4 U6787 ( .INP(n5874), .Z(n5963) );
  NBUFFX4 U6788 ( .INP(n5874), .Z(n5964) );
  INVX0 U6789 ( .INP(wraddr[1]), .ZN(n7363) );
  INVX0 U6790 ( .INP(wraddr[3]), .ZN(n7365) );
  NOR2X0 U6791 ( .IN1(n7364), .IN2(wraddr[3]), .QN(n389) );
  NOR2X0 U6792 ( .IN1(wraddr[2]), .IN2(wraddr[3]), .QN(n394) );
  NOR2X0 U6793 ( .IN1(n7362), .IN2(wraddr[1]), .QN(n380) );
  NOR2X0 U6794 ( .IN1(wraddr[0]), .IN2(wraddr[1]), .QN(n382) );
  INVX0 U6795 ( .INP(wraddr[2]), .ZN(n7364) );
  INVX0 U6796 ( .INP(wraddr[0]), .ZN(n7362) );
  AND4X4 U6797 ( .IN1(wraddr[5]), .IN2(wraddr[4]), .IN3(n270), .IN4(n7368), 
        .Q(n323) );
  AND4X4 U6798 ( .IN1(wraddr[6]), .IN2(wraddr[4]), .IN3(n270), .IN4(n7367), 
        .Q(n289) );
  NOR2X0 U6799 ( .IN1(wraddr[7]), .IN2(n8), .QN(n270) );
  AND4X4 U6800 ( .IN1(n7368), .IN2(n7366), .IN3(n7367), .IN4(n270), .Q(n374)
         );
  AND4X4 U6801 ( .IN1(wraddr[6]), .IN2(wraddr[5]), .IN3(n270), .IN4(n7366), 
        .Q(n272) );
  AND4X4 U6802 ( .IN1(wraddr[6]), .IN2(wraddr[5]), .IN3(wraddr[4]), .IN4(n270), 
        .Q(n239) );
  INVX0 U6803 ( .INP(n52), .ZN(n5976) );
  INVX0 U6804 ( .INP(n52), .ZN(n5977) );
  INVX0 U6805 ( .INP(n52), .ZN(n5978) );
  INVX0 U6806 ( .INP(n397), .ZN(n5982) );
  INVX0 U6807 ( .INP(n397), .ZN(n5983) );
  INVX0 U6808 ( .INP(n397), .ZN(n5984) );
  INVX0 U6809 ( .INP(n396), .ZN(n5988) );
  INVX0 U6810 ( .INP(n396), .ZN(n5989) );
  INVX0 U6811 ( .INP(n396), .ZN(n5990) );
  INVX0 U6812 ( .INP(n395), .ZN(n5994) );
  INVX0 U6813 ( .INP(n395), .ZN(n5995) );
  INVX0 U6814 ( .INP(n395), .ZN(n5996) );
  INVX0 U6815 ( .INP(n393), .ZN(n6000) );
  INVX0 U6816 ( .INP(n393), .ZN(n6001) );
  INVX0 U6817 ( .INP(n393), .ZN(n6002) );
  INVX0 U6818 ( .INP(n392), .ZN(n6006) );
  INVX0 U6819 ( .INP(n392), .ZN(n6007) );
  INVX0 U6820 ( .INP(n392), .ZN(n6008) );
  INVX0 U6821 ( .INP(n391), .ZN(n6012) );
  INVX0 U6822 ( .INP(n391), .ZN(n6013) );
  INVX0 U6823 ( .INP(n391), .ZN(n6014) );
  INVX0 U6824 ( .INP(n390), .ZN(n6018) );
  INVX0 U6825 ( .INP(n390), .ZN(n6019) );
  INVX0 U6826 ( .INP(n390), .ZN(n6020) );
  INVX0 U6827 ( .INP(n388), .ZN(n6024) );
  INVX0 U6828 ( .INP(n388), .ZN(n6025) );
  INVX0 U6829 ( .INP(n388), .ZN(n6026) );
  INVX0 U6830 ( .INP(n387), .ZN(n6030) );
  INVX0 U6831 ( .INP(n387), .ZN(n6031) );
  INVX0 U6832 ( .INP(n387), .ZN(n6032) );
  INVX0 U6833 ( .INP(n386), .ZN(n6036) );
  INVX0 U6834 ( .INP(n386), .ZN(n6037) );
  INVX0 U6835 ( .INP(n386), .ZN(n6038) );
  INVX0 U6836 ( .INP(n385), .ZN(n6042) );
  INVX0 U6837 ( .INP(n385), .ZN(n6043) );
  INVX0 U6838 ( .INP(n385), .ZN(n6044) );
  INVX0 U6839 ( .INP(n383), .ZN(n6048) );
  INVX0 U6840 ( .INP(n383), .ZN(n6049) );
  INVX0 U6841 ( .INP(n383), .ZN(n6050) );
  INVX0 U6842 ( .INP(n381), .ZN(n6054) );
  INVX0 U6843 ( .INP(n381), .ZN(n6055) );
  INVX0 U6844 ( .INP(n381), .ZN(n6056) );
  INVX0 U6845 ( .INP(n379), .ZN(n6060) );
  INVX0 U6846 ( .INP(n379), .ZN(n6061) );
  INVX0 U6847 ( .INP(n379), .ZN(n6062) );
  INVX0 U6848 ( .INP(n377), .ZN(n6066) );
  INVX0 U6849 ( .INP(n377), .ZN(n6067) );
  INVX0 U6850 ( .INP(n377), .ZN(n6068) );
  INVX0 U6851 ( .INP(n373), .ZN(n6072) );
  INVX0 U6852 ( .INP(n373), .ZN(n6073) );
  INVX0 U6853 ( .INP(n373), .ZN(n6074) );
  INVX0 U6854 ( .INP(n372), .ZN(n6078) );
  INVX0 U6855 ( .INP(n372), .ZN(n6079) );
  INVX0 U6856 ( .INP(n372), .ZN(n6080) );
  INVX0 U6857 ( .INP(n371), .ZN(n6084) );
  INVX0 U6858 ( .INP(n371), .ZN(n6085) );
  INVX0 U6859 ( .INP(n371), .ZN(n6086) );
  INVX0 U6860 ( .INP(n370), .ZN(n6090) );
  INVX0 U6861 ( .INP(n370), .ZN(n6091) );
  INVX0 U6862 ( .INP(n370), .ZN(n6092) );
  INVX0 U6863 ( .INP(n369), .ZN(n6096) );
  INVX0 U6864 ( .INP(n369), .ZN(n6097) );
  INVX0 U6865 ( .INP(n369), .ZN(n6098) );
  INVX0 U6866 ( .INP(n368), .ZN(n6102) );
  INVX0 U6867 ( .INP(n368), .ZN(n6103) );
  INVX0 U6868 ( .INP(n368), .ZN(n6104) );
  INVX0 U6869 ( .INP(n367), .ZN(n6108) );
  INVX0 U6870 ( .INP(n367), .ZN(n6109) );
  INVX0 U6871 ( .INP(n367), .ZN(n6110) );
  INVX0 U6872 ( .INP(n366), .ZN(n6114) );
  INVX0 U6873 ( .INP(n366), .ZN(n6115) );
  INVX0 U6874 ( .INP(n366), .ZN(n6116) );
  INVX0 U6875 ( .INP(n365), .ZN(n6120) );
  INVX0 U6876 ( .INP(n365), .ZN(n6121) );
  INVX0 U6877 ( .INP(n365), .ZN(n6122) );
  INVX0 U6878 ( .INP(n364), .ZN(n6126) );
  INVX0 U6879 ( .INP(n364), .ZN(n6127) );
  INVX0 U6880 ( .INP(n364), .ZN(n6128) );
  INVX0 U6881 ( .INP(n363), .ZN(n6132) );
  INVX0 U6882 ( .INP(n363), .ZN(n6133) );
  INVX0 U6883 ( .INP(n363), .ZN(n6134) );
  INVX0 U6884 ( .INP(n362), .ZN(n6138) );
  INVX0 U6885 ( .INP(n362), .ZN(n6139) );
  INVX0 U6886 ( .INP(n362), .ZN(n6140) );
  INVX0 U6887 ( .INP(n361), .ZN(n6144) );
  INVX0 U6888 ( .INP(n361), .ZN(n6145) );
  INVX0 U6889 ( .INP(n361), .ZN(n6146) );
  INVX0 U6890 ( .INP(n360), .ZN(n6150) );
  INVX0 U6891 ( .INP(n360), .ZN(n6151) );
  INVX0 U6892 ( .INP(n360), .ZN(n6152) );
  INVX0 U6893 ( .INP(n359), .ZN(n6156) );
  INVX0 U6894 ( .INP(n359), .ZN(n6157) );
  INVX0 U6895 ( .INP(n359), .ZN(n6158) );
  INVX0 U6896 ( .INP(n358), .ZN(n6162) );
  INVX0 U6897 ( .INP(n358), .ZN(n6163) );
  INVX0 U6898 ( .INP(n358), .ZN(n6164) );
  INVX0 U6899 ( .INP(n356), .ZN(n6168) );
  INVX0 U6900 ( .INP(n356), .ZN(n6169) );
  INVX0 U6901 ( .INP(n356), .ZN(n6170) );
  INVX0 U6902 ( .INP(n355), .ZN(n6174) );
  INVX0 U6903 ( .INP(n355), .ZN(n6175) );
  INVX0 U6904 ( .INP(n355), .ZN(n6176) );
  INVX0 U6905 ( .INP(n354), .ZN(n6180) );
  INVX0 U6906 ( .INP(n354), .ZN(n6181) );
  INVX0 U6907 ( .INP(n354), .ZN(n6182) );
  INVX0 U6908 ( .INP(n353), .ZN(n6186) );
  INVX0 U6909 ( .INP(n353), .ZN(n6187) );
  INVX0 U6910 ( .INP(n353), .ZN(n6188) );
  INVX0 U6911 ( .INP(n352), .ZN(n6192) );
  INVX0 U6912 ( .INP(n352), .ZN(n6193) );
  INVX0 U6913 ( .INP(n352), .ZN(n6194) );
  INVX0 U6914 ( .INP(n351), .ZN(n6198) );
  INVX0 U6915 ( .INP(n351), .ZN(n6199) );
  INVX0 U6916 ( .INP(n351), .ZN(n6200) );
  INVX0 U6917 ( .INP(n350), .ZN(n6204) );
  INVX0 U6918 ( .INP(n350), .ZN(n6205) );
  INVX0 U6919 ( .INP(n350), .ZN(n6206) );
  INVX0 U6920 ( .INP(n349), .ZN(n6210) );
  INVX0 U6921 ( .INP(n349), .ZN(n6211) );
  INVX0 U6922 ( .INP(n349), .ZN(n6212) );
  INVX0 U6923 ( .INP(n348), .ZN(n6216) );
  INVX0 U6924 ( .INP(n348), .ZN(n6217) );
  INVX0 U6925 ( .INP(n348), .ZN(n6218) );
  INVX0 U6926 ( .INP(n347), .ZN(n6222) );
  INVX0 U6927 ( .INP(n347), .ZN(n6223) );
  INVX0 U6928 ( .INP(n347), .ZN(n6224) );
  INVX0 U6929 ( .INP(n346), .ZN(n6228) );
  INVX0 U6930 ( .INP(n346), .ZN(n6229) );
  INVX0 U6931 ( .INP(n346), .ZN(n6230) );
  INVX0 U6932 ( .INP(n345), .ZN(n6234) );
  INVX0 U6933 ( .INP(n345), .ZN(n6235) );
  INVX0 U6934 ( .INP(n345), .ZN(n6236) );
  INVX0 U6935 ( .INP(n344), .ZN(n6240) );
  INVX0 U6936 ( .INP(n344), .ZN(n6241) );
  INVX0 U6937 ( .INP(n344), .ZN(n6242) );
  INVX0 U6938 ( .INP(n343), .ZN(n6246) );
  INVX0 U6939 ( .INP(n343), .ZN(n6247) );
  INVX0 U6940 ( .INP(n343), .ZN(n6248) );
  INVX0 U6941 ( .INP(n342), .ZN(n6252) );
  INVX0 U6942 ( .INP(n342), .ZN(n6253) );
  INVX0 U6943 ( .INP(n342), .ZN(n6254) );
  INVX0 U6944 ( .INP(n341), .ZN(n6258) );
  INVX0 U6945 ( .INP(n341), .ZN(n6259) );
  INVX0 U6946 ( .INP(n341), .ZN(n6260) );
  INVX0 U6947 ( .INP(n339), .ZN(n6264) );
  INVX0 U6948 ( .INP(n339), .ZN(n6265) );
  INVX0 U6949 ( .INP(n339), .ZN(n6266) );
  INVX0 U6950 ( .INP(n338), .ZN(n6270) );
  INVX0 U6951 ( .INP(n338), .ZN(n6271) );
  INVX0 U6952 ( .INP(n338), .ZN(n6272) );
  INVX0 U6953 ( .INP(n337), .ZN(n6276) );
  INVX0 U6954 ( .INP(n337), .ZN(n6277) );
  INVX0 U6955 ( .INP(n337), .ZN(n6278) );
  INVX0 U6956 ( .INP(n336), .ZN(n6282) );
  INVX0 U6957 ( .INP(n336), .ZN(n6283) );
  INVX0 U6958 ( .INP(n336), .ZN(n6284) );
  INVX0 U6959 ( .INP(n335), .ZN(n6288) );
  INVX0 U6960 ( .INP(n335), .ZN(n6289) );
  INVX0 U6961 ( .INP(n335), .ZN(n6290) );
  INVX0 U6962 ( .INP(n334), .ZN(n6294) );
  INVX0 U6963 ( .INP(n334), .ZN(n6295) );
  INVX0 U6964 ( .INP(n334), .ZN(n6296) );
  INVX0 U6965 ( .INP(n333), .ZN(n6300) );
  INVX0 U6966 ( .INP(n333), .ZN(n6301) );
  INVX0 U6967 ( .INP(n333), .ZN(n6302) );
  INVX0 U6968 ( .INP(n332), .ZN(n6306) );
  INVX0 U6969 ( .INP(n332), .ZN(n6307) );
  INVX0 U6970 ( .INP(n332), .ZN(n6308) );
  INVX0 U6971 ( .INP(n331), .ZN(n6312) );
  INVX0 U6972 ( .INP(n331), .ZN(n6313) );
  INVX0 U6973 ( .INP(n331), .ZN(n6314) );
  INVX0 U6974 ( .INP(n330), .ZN(n6318) );
  INVX0 U6975 ( .INP(n330), .ZN(n6319) );
  INVX0 U6976 ( .INP(n330), .ZN(n6320) );
  INVX0 U6977 ( .INP(n329), .ZN(n6324) );
  INVX0 U6978 ( .INP(n329), .ZN(n6325) );
  INVX0 U6979 ( .INP(n329), .ZN(n6326) );
  INVX0 U6980 ( .INP(n328), .ZN(n6330) );
  INVX0 U6981 ( .INP(n328), .ZN(n6331) );
  INVX0 U6982 ( .INP(n328), .ZN(n6332) );
  INVX0 U6983 ( .INP(n327), .ZN(n6336) );
  INVX0 U6984 ( .INP(n327), .ZN(n6337) );
  INVX0 U6985 ( .INP(n327), .ZN(n6338) );
  INVX0 U6986 ( .INP(n326), .ZN(n6342) );
  INVX0 U6987 ( .INP(n326), .ZN(n6343) );
  INVX0 U6988 ( .INP(n326), .ZN(n6344) );
  INVX0 U6989 ( .INP(n325), .ZN(n6348) );
  INVX0 U6990 ( .INP(n325), .ZN(n6349) );
  INVX0 U6991 ( .INP(n325), .ZN(n6350) );
  INVX0 U6992 ( .INP(n324), .ZN(n6354) );
  INVX0 U6993 ( .INP(n324), .ZN(n6355) );
  INVX0 U6994 ( .INP(n324), .ZN(n6356) );
  INVX0 U6995 ( .INP(n322), .ZN(n6360) );
  INVX0 U6996 ( .INP(n322), .ZN(n6361) );
  INVX0 U6997 ( .INP(n322), .ZN(n6362) );
  INVX0 U6998 ( .INP(n321), .ZN(n6366) );
  INVX0 U6999 ( .INP(n321), .ZN(n6367) );
  INVX0 U7000 ( .INP(n321), .ZN(n6368) );
  INVX0 U7001 ( .INP(n320), .ZN(n6372) );
  INVX0 U7002 ( .INP(n320), .ZN(n6373) );
  INVX0 U7003 ( .INP(n320), .ZN(n6374) );
  INVX0 U7004 ( .INP(n319), .ZN(n6378) );
  INVX0 U7005 ( .INP(n319), .ZN(n6379) );
  INVX0 U7006 ( .INP(n319), .ZN(n6380) );
  INVX0 U7007 ( .INP(n318), .ZN(n6384) );
  INVX0 U7008 ( .INP(n318), .ZN(n6385) );
  INVX0 U7009 ( .INP(n318), .ZN(n6386) );
  INVX0 U7010 ( .INP(n317), .ZN(n6390) );
  INVX0 U7011 ( .INP(n317), .ZN(n6391) );
  INVX0 U7012 ( .INP(n317), .ZN(n6392) );
  INVX0 U7013 ( .INP(n316), .ZN(n6396) );
  INVX0 U7014 ( .INP(n316), .ZN(n6397) );
  INVX0 U7015 ( .INP(n316), .ZN(n6398) );
  INVX0 U7016 ( .INP(n315), .ZN(n6402) );
  INVX0 U7017 ( .INP(n315), .ZN(n6403) );
  INVX0 U7018 ( .INP(n315), .ZN(n6404) );
  INVX0 U7019 ( .INP(n314), .ZN(n6408) );
  INVX0 U7020 ( .INP(n314), .ZN(n6409) );
  INVX0 U7021 ( .INP(n314), .ZN(n6410) );
  INVX0 U7022 ( .INP(n313), .ZN(n6414) );
  INVX0 U7023 ( .INP(n313), .ZN(n6415) );
  INVX0 U7024 ( .INP(n313), .ZN(n6416) );
  INVX0 U7025 ( .INP(n312), .ZN(n6420) );
  INVX0 U7026 ( .INP(n312), .ZN(n6421) );
  INVX0 U7027 ( .INP(n312), .ZN(n6422) );
  INVX0 U7028 ( .INP(n311), .ZN(n6426) );
  INVX0 U7029 ( .INP(n311), .ZN(n6427) );
  INVX0 U7030 ( .INP(n311), .ZN(n6428) );
  INVX0 U7031 ( .INP(n310), .ZN(n6432) );
  INVX0 U7032 ( .INP(n310), .ZN(n6433) );
  INVX0 U7033 ( .INP(n310), .ZN(n6434) );
  INVX0 U7034 ( .INP(n309), .ZN(n6438) );
  INVX0 U7035 ( .INP(n309), .ZN(n6439) );
  INVX0 U7036 ( .INP(n309), .ZN(n6440) );
  INVX0 U7037 ( .INP(n308), .ZN(n6444) );
  INVX0 U7038 ( .INP(n308), .ZN(n6445) );
  INVX0 U7039 ( .INP(n308), .ZN(n6446) );
  INVX0 U7040 ( .INP(n307), .ZN(n6450) );
  INVX0 U7041 ( .INP(n307), .ZN(n6451) );
  INVX0 U7042 ( .INP(n307), .ZN(n6452) );
  INVX0 U7043 ( .INP(n305), .ZN(n6456) );
  INVX0 U7044 ( .INP(n305), .ZN(n6457) );
  INVX0 U7045 ( .INP(n305), .ZN(n6458) );
  INVX0 U7046 ( .INP(n304), .ZN(n6462) );
  INVX0 U7047 ( .INP(n304), .ZN(n6463) );
  INVX0 U7048 ( .INP(n304), .ZN(n6464) );
  INVX0 U7049 ( .INP(n303), .ZN(n6468) );
  INVX0 U7050 ( .INP(n303), .ZN(n6469) );
  INVX0 U7051 ( .INP(n303), .ZN(n6470) );
  INVX0 U7052 ( .INP(n302), .ZN(n6474) );
  INVX0 U7053 ( .INP(n302), .ZN(n6475) );
  INVX0 U7054 ( .INP(n302), .ZN(n6476) );
  INVX0 U7055 ( .INP(n301), .ZN(n6480) );
  INVX0 U7056 ( .INP(n301), .ZN(n6481) );
  INVX0 U7057 ( .INP(n301), .ZN(n6482) );
  INVX0 U7058 ( .INP(n300), .ZN(n6486) );
  INVX0 U7059 ( .INP(n300), .ZN(n6487) );
  INVX0 U7060 ( .INP(n300), .ZN(n6488) );
  INVX0 U7061 ( .INP(n299), .ZN(n6492) );
  INVX0 U7062 ( .INP(n299), .ZN(n6493) );
  INVX0 U7063 ( .INP(n299), .ZN(n6494) );
  INVX0 U7064 ( .INP(n298), .ZN(n6498) );
  INVX0 U7065 ( .INP(n298), .ZN(n6499) );
  INVX0 U7066 ( .INP(n298), .ZN(n6500) );
  INVX0 U7067 ( .INP(n297), .ZN(n6504) );
  INVX0 U7068 ( .INP(n297), .ZN(n6505) );
  INVX0 U7069 ( .INP(n297), .ZN(n6506) );
  INVX0 U7070 ( .INP(n296), .ZN(n6510) );
  INVX0 U7071 ( .INP(n296), .ZN(n6511) );
  INVX0 U7072 ( .INP(n296), .ZN(n6512) );
  INVX0 U7073 ( .INP(n295), .ZN(n6516) );
  INVX0 U7074 ( .INP(n295), .ZN(n6517) );
  INVX0 U7075 ( .INP(n295), .ZN(n6518) );
  INVX0 U7076 ( .INP(n294), .ZN(n6522) );
  INVX0 U7077 ( .INP(n294), .ZN(n6523) );
  INVX0 U7078 ( .INP(n294), .ZN(n6524) );
  INVX0 U7079 ( .INP(n293), .ZN(n6528) );
  INVX0 U7080 ( .INP(n293), .ZN(n6529) );
  INVX0 U7081 ( .INP(n293), .ZN(n6530) );
  INVX0 U7082 ( .INP(n292), .ZN(n6534) );
  INVX0 U7083 ( .INP(n292), .ZN(n6535) );
  INVX0 U7084 ( .INP(n292), .ZN(n6536) );
  INVX0 U7085 ( .INP(n291), .ZN(n6540) );
  INVX0 U7086 ( .INP(n291), .ZN(n6541) );
  INVX0 U7087 ( .INP(n291), .ZN(n6542) );
  INVX0 U7088 ( .INP(n290), .ZN(n6546) );
  INVX0 U7089 ( .INP(n290), .ZN(n6547) );
  INVX0 U7090 ( .INP(n290), .ZN(n6548) );
  INVX0 U7091 ( .INP(n288), .ZN(n6552) );
  INVX0 U7092 ( .INP(n288), .ZN(n6553) );
  INVX0 U7093 ( .INP(n288), .ZN(n6554) );
  INVX0 U7094 ( .INP(n287), .ZN(n6558) );
  INVX0 U7095 ( .INP(n287), .ZN(n6559) );
  INVX0 U7096 ( .INP(n287), .ZN(n6560) );
  INVX0 U7097 ( .INP(n286), .ZN(n6564) );
  INVX0 U7098 ( .INP(n286), .ZN(n6565) );
  INVX0 U7099 ( .INP(n286), .ZN(n6566) );
  INVX0 U7100 ( .INP(n285), .ZN(n6570) );
  INVX0 U7101 ( .INP(n285), .ZN(n6571) );
  INVX0 U7102 ( .INP(n285), .ZN(n6572) );
  INVX0 U7103 ( .INP(n284), .ZN(n6576) );
  INVX0 U7104 ( .INP(n284), .ZN(n6577) );
  INVX0 U7105 ( .INP(n284), .ZN(n6578) );
  INVX0 U7106 ( .INP(n283), .ZN(n6582) );
  INVX0 U7107 ( .INP(n283), .ZN(n6583) );
  INVX0 U7108 ( .INP(n283), .ZN(n6584) );
  INVX0 U7109 ( .INP(n282), .ZN(n6588) );
  INVX0 U7110 ( .INP(n282), .ZN(n6589) );
  INVX0 U7111 ( .INP(n282), .ZN(n6590) );
  INVX0 U7112 ( .INP(n281), .ZN(n6594) );
  INVX0 U7113 ( .INP(n281), .ZN(n6595) );
  INVX0 U7114 ( .INP(n281), .ZN(n6596) );
  INVX0 U7115 ( .INP(n280), .ZN(n6600) );
  INVX0 U7116 ( .INP(n280), .ZN(n6601) );
  INVX0 U7117 ( .INP(n280), .ZN(n6602) );
  INVX0 U7118 ( .INP(n279), .ZN(n6606) );
  INVX0 U7119 ( .INP(n279), .ZN(n6607) );
  INVX0 U7120 ( .INP(n279), .ZN(n6608) );
  INVX0 U7121 ( .INP(n278), .ZN(n6612) );
  INVX0 U7122 ( .INP(n278), .ZN(n6613) );
  INVX0 U7123 ( .INP(n278), .ZN(n6614) );
  INVX0 U7124 ( .INP(n277), .ZN(n6618) );
  INVX0 U7125 ( .INP(n277), .ZN(n6619) );
  INVX0 U7126 ( .INP(n277), .ZN(n6620) );
  INVX0 U7127 ( .INP(n276), .ZN(n6624) );
  INVX0 U7128 ( .INP(n276), .ZN(n6625) );
  INVX0 U7129 ( .INP(n276), .ZN(n6626) );
  INVX0 U7130 ( .INP(n275), .ZN(n6630) );
  INVX0 U7131 ( .INP(n275), .ZN(n6631) );
  INVX0 U7132 ( .INP(n275), .ZN(n6632) );
  INVX0 U7133 ( .INP(n274), .ZN(n6636) );
  INVX0 U7134 ( .INP(n274), .ZN(n6637) );
  INVX0 U7135 ( .INP(n274), .ZN(n6638) );
  INVX0 U7136 ( .INP(n273), .ZN(n6642) );
  INVX0 U7137 ( .INP(n273), .ZN(n6643) );
  INVX0 U7138 ( .INP(n273), .ZN(n6644) );
  INVX0 U7139 ( .INP(n271), .ZN(n6648) );
  INVX0 U7140 ( .INP(n271), .ZN(n6649) );
  INVX0 U7141 ( .INP(n271), .ZN(n6650) );
  INVX0 U7142 ( .INP(n268), .ZN(n6654) );
  INVX0 U7143 ( .INP(n268), .ZN(n6655) );
  INVX0 U7144 ( .INP(n268), .ZN(n6656) );
  INVX0 U7145 ( .INP(n266), .ZN(n6660) );
  INVX0 U7146 ( .INP(n266), .ZN(n6661) );
  INVX0 U7147 ( .INP(n266), .ZN(n6662) );
  INVX0 U7148 ( .INP(n264), .ZN(n6666) );
  INVX0 U7149 ( .INP(n264), .ZN(n6667) );
  INVX0 U7150 ( .INP(n264), .ZN(n6668) );
  INVX0 U7151 ( .INP(n262), .ZN(n6672) );
  INVX0 U7152 ( .INP(n262), .ZN(n6673) );
  INVX0 U7153 ( .INP(n262), .ZN(n6674) );
  INVX0 U7154 ( .INP(n260), .ZN(n6678) );
  INVX0 U7155 ( .INP(n260), .ZN(n6679) );
  INVX0 U7156 ( .INP(n260), .ZN(n6680) );
  INVX0 U7157 ( .INP(n258), .ZN(n6684) );
  INVX0 U7158 ( .INP(n258), .ZN(n6685) );
  INVX0 U7159 ( .INP(n258), .ZN(n6686) );
  INVX0 U7160 ( .INP(n256), .ZN(n6690) );
  INVX0 U7161 ( .INP(n256), .ZN(n6691) );
  INVX0 U7162 ( .INP(n256), .ZN(n6692) );
  INVX0 U7163 ( .INP(n254), .ZN(n6696) );
  INVX0 U7164 ( .INP(n254), .ZN(n6697) );
  INVX0 U7165 ( .INP(n254), .ZN(n6698) );
  INVX0 U7166 ( .INP(n252), .ZN(n6702) );
  INVX0 U7167 ( .INP(n252), .ZN(n6703) );
  INVX0 U7168 ( .INP(n252), .ZN(n6704) );
  INVX0 U7169 ( .INP(n250), .ZN(n6708) );
  INVX0 U7170 ( .INP(n250), .ZN(n6709) );
  INVX0 U7171 ( .INP(n250), .ZN(n6710) );
  INVX0 U7172 ( .INP(n248), .ZN(n6714) );
  INVX0 U7173 ( .INP(n248), .ZN(n6715) );
  INVX0 U7174 ( .INP(n248), .ZN(n6716) );
  INVX0 U7175 ( .INP(n246), .ZN(n6720) );
  INVX0 U7176 ( .INP(n246), .ZN(n6721) );
  INVX0 U7177 ( .INP(n246), .ZN(n6722) );
  INVX0 U7178 ( .INP(n244), .ZN(n6726) );
  INVX0 U7179 ( .INP(n244), .ZN(n6727) );
  INVX0 U7180 ( .INP(n244), .ZN(n6728) );
  INVX0 U7181 ( .INP(n242), .ZN(n6732) );
  INVX0 U7182 ( .INP(n242), .ZN(n6733) );
  INVX0 U7183 ( .INP(n242), .ZN(n6734) );
  INVX0 U7184 ( .INP(n240), .ZN(n6738) );
  INVX0 U7185 ( .INP(n240), .ZN(n6739) );
  INVX0 U7186 ( .INP(n240), .ZN(n6740) );
  INVX0 U7187 ( .INP(n206), .ZN(n7085) );
  INVX0 U7188 ( .INP(n206), .ZN(n7086) );
  INVX0 U7189 ( .INP(n206), .ZN(n7087) );
  INVX0 U7190 ( .INP(n7102), .ZN(n7099) );
  INVX0 U7191 ( .INP(n7101), .ZN(n7100) );
  INVX0 U7192 ( .INP(n7339), .ZN(n7104) );
  INVX0 U7193 ( .INP(n7340), .ZN(n7105) );
  INVX0 U7194 ( .INP(n7348), .ZN(n7106) );
  INVX0 U7195 ( .INP(n7338), .ZN(n7107) );
  INVX0 U7196 ( .INP(n7339), .ZN(n7108) );
  INVX0 U7197 ( .INP(n7341), .ZN(n7109) );
  INVX0 U7198 ( .INP(n7342), .ZN(n7110) );
  INVX0 U7199 ( .INP(n7343), .ZN(n7111) );
  INVX0 U7200 ( .INP(n7347), .ZN(n7112) );
  INVX0 U7201 ( .INP(n7336), .ZN(n7113) );
  INVX0 U7202 ( .INP(n7337), .ZN(n7114) );
  INVX0 U7203 ( .INP(n7338), .ZN(n7115) );
  INVX0 U7204 ( .INP(n7339), .ZN(n7116) );
  INVX0 U7205 ( .INP(n7341), .ZN(n7117) );
  INVX0 U7206 ( .INP(n7342), .ZN(n7118) );
  INVX0 U7207 ( .INP(n7348), .ZN(n7119) );
  INVX0 U7208 ( .INP(n7349), .ZN(n7120) );
  INVX0 U7209 ( .INP(n7350), .ZN(n7121) );
  INVX0 U7210 ( .INP(n7351), .ZN(n7122) );
  INVX0 U7211 ( .INP(n7352), .ZN(n7123) );
  INVX0 U7212 ( .INP(n7344), .ZN(n7124) );
  INVX0 U7213 ( .INP(n7343), .ZN(n7125) );
  INVX0 U7214 ( .INP(n7334), .ZN(n7126) );
  INVX0 U7215 ( .INP(n7353), .ZN(n7127) );
  INVX0 U7216 ( .INP(n7335), .ZN(n7128) );
  INVX0 U7217 ( .INP(n7352), .ZN(n7129) );
  INVX0 U7218 ( .INP(n7337), .ZN(n7130) );
  INVX0 U7219 ( .INP(n7352), .ZN(n7131) );
  INVX0 U7220 ( .INP(n7352), .ZN(n7132) );
  INVX0 U7221 ( .INP(n7352), .ZN(n7133) );
  INVX0 U7222 ( .INP(n7352), .ZN(n7134) );
  INVX0 U7223 ( .INP(n7352), .ZN(n7135) );
  INVX0 U7224 ( .INP(n7352), .ZN(n7136) );
  INVX0 U7225 ( .INP(n7351), .ZN(n7137) );
  INVX0 U7226 ( .INP(n7351), .ZN(n7138) );
  INVX0 U7227 ( .INP(n7351), .ZN(n7139) );
  INVX0 U7228 ( .INP(n7351), .ZN(n7140) );
  INVX0 U7229 ( .INP(n7351), .ZN(n7141) );
  INVX0 U7230 ( .INP(n7351), .ZN(n7142) );
  INVX0 U7231 ( .INP(n7350), .ZN(n7143) );
  INVX0 U7232 ( .INP(n7350), .ZN(n7144) );
  INVX0 U7233 ( .INP(n7350), .ZN(n7145) );
  INVX0 U7234 ( .INP(n7350), .ZN(n7146) );
  INVX0 U7235 ( .INP(n7350), .ZN(n7147) );
  INVX0 U7236 ( .INP(n7350), .ZN(n7148) );
  INVX0 U7237 ( .INP(n7349), .ZN(n7149) );
  INVX0 U7238 ( .INP(n7349), .ZN(n7150) );
  INVX0 U7239 ( .INP(n7349), .ZN(n7151) );
  INVX0 U7240 ( .INP(n7349), .ZN(n7152) );
  INVX0 U7241 ( .INP(n7349), .ZN(n7153) );
  INVX0 U7242 ( .INP(n7349), .ZN(n7154) );
  INVX0 U7243 ( .INP(n7348), .ZN(n7155) );
  INVX0 U7244 ( .INP(n7348), .ZN(n7156) );
  INVX0 U7245 ( .INP(n7348), .ZN(n7157) );
  INVX0 U7246 ( .INP(n7348), .ZN(n7158) );
  INVX0 U7247 ( .INP(n7348), .ZN(n7159) );
  INVX0 U7248 ( .INP(n7348), .ZN(n7160) );
  INVX0 U7249 ( .INP(n7347), .ZN(n7161) );
  INVX0 U7250 ( .INP(n7347), .ZN(n7162) );
  INVX0 U7251 ( .INP(n7347), .ZN(n7163) );
  INVX0 U7252 ( .INP(n7347), .ZN(n7164) );
  INVX0 U7253 ( .INP(n7347), .ZN(n7165) );
  INVX0 U7254 ( .INP(n7347), .ZN(n7166) );
  INVX0 U7255 ( .INP(n7346), .ZN(n7167) );
  INVX0 U7256 ( .INP(n7346), .ZN(n7168) );
  INVX0 U7257 ( .INP(n7346), .ZN(n7169) );
  INVX0 U7258 ( .INP(n7346), .ZN(n7170) );
  INVX0 U7259 ( .INP(n7346), .ZN(n7171) );
  INVX0 U7260 ( .INP(n7346), .ZN(n7172) );
  INVX0 U7261 ( .INP(n7345), .ZN(n7173) );
  INVX0 U7262 ( .INP(n7345), .ZN(n7174) );
  INVX0 U7263 ( .INP(n7345), .ZN(n7175) );
  INVX0 U7264 ( .INP(n7345), .ZN(n7176) );
  INVX0 U7265 ( .INP(n7345), .ZN(n7177) );
  INVX0 U7266 ( .INP(n7345), .ZN(n7178) );
  INVX0 U7267 ( .INP(n7344), .ZN(n7179) );
  INVX0 U7268 ( .INP(n7344), .ZN(n7180) );
  INVX0 U7269 ( .INP(n7344), .ZN(n7181) );
  INVX0 U7270 ( .INP(n7344), .ZN(n7182) );
  INVX0 U7271 ( .INP(n7344), .ZN(n7183) );
  INVX0 U7272 ( .INP(n7344), .ZN(n7184) );
  INVX0 U7273 ( .INP(n7343), .ZN(n7185) );
  INVX0 U7274 ( .INP(n7343), .ZN(n7186) );
  INVX0 U7275 ( .INP(n7343), .ZN(n7187) );
  INVX0 U7276 ( .INP(n7343), .ZN(n7188) );
  INVX0 U7277 ( .INP(n7343), .ZN(n7189) );
  INVX0 U7278 ( .INP(n7343), .ZN(n7190) );
  INVX0 U7279 ( .INP(n7342), .ZN(n7191) );
  INVX0 U7280 ( .INP(n7342), .ZN(n7192) );
  INVX0 U7281 ( .INP(n7342), .ZN(n7193) );
  INVX0 U7282 ( .INP(n7342), .ZN(n7194) );
  INVX0 U7283 ( .INP(n7342), .ZN(n7195) );
  INVX0 U7284 ( .INP(n7342), .ZN(n7196) );
  INVX0 U7285 ( .INP(n7341), .ZN(n7197) );
  INVX0 U7286 ( .INP(n7341), .ZN(n7198) );
  INVX0 U7287 ( .INP(n7341), .ZN(n7199) );
  INVX0 U7288 ( .INP(n7341), .ZN(n7200) );
  INVX0 U7289 ( .INP(n7341), .ZN(n7201) );
  INVX0 U7290 ( .INP(n7341), .ZN(n7202) );
  INVX0 U7291 ( .INP(n7340), .ZN(n7203) );
  INVX0 U7292 ( .INP(n7340), .ZN(n7204) );
  INVX0 U7293 ( .INP(n7340), .ZN(n7205) );
  INVX0 U7294 ( .INP(n7340), .ZN(n7206) );
  INVX0 U7295 ( .INP(n7340), .ZN(n7207) );
  INVX0 U7296 ( .INP(n7340), .ZN(n7208) );
  INVX0 U7297 ( .INP(n7335), .ZN(n7209) );
  INVX0 U7298 ( .INP(n7336), .ZN(n7210) );
  INVX0 U7299 ( .INP(n7358), .ZN(n7211) );
  INVX0 U7300 ( .INP(n7355), .ZN(n7212) );
  INVX0 U7301 ( .INP(n7354), .ZN(n7213) );
  INVX0 U7302 ( .INP(n7345), .ZN(n7214) );
  INVX0 U7303 ( .INP(n7356), .ZN(n7215) );
  INVX0 U7304 ( .INP(n7344), .ZN(n7216) );
  INVX0 U7305 ( .INP(n7347), .ZN(n7217) );
  INVX0 U7306 ( .INP(n7352), .ZN(n7218) );
  INVX0 U7307 ( .INP(n7353), .ZN(n7219) );
  INVX0 U7308 ( .INP(n7339), .ZN(n7220) );
  INVX0 U7309 ( .INP(n7353), .ZN(n7221) );
  INVX0 U7310 ( .INP(n7335), .ZN(n7222) );
  INVX0 U7311 ( .INP(n7358), .ZN(n7223) );
  INVX0 U7312 ( .INP(n7348), .ZN(n7224) );
  INVX0 U7313 ( .INP(n7340), .ZN(n7225) );
  INVX0 U7314 ( .INP(n7349), .ZN(n7226) );
  INVX0 U7315 ( .INP(n7346), .ZN(n7227) );
  INVX0 U7316 ( .INP(n7358), .ZN(n7228) );
  INVX0 U7317 ( .INP(n7354), .ZN(n7229) );
  INVX0 U7318 ( .INP(n7355), .ZN(n7230) );
  INVX0 U7319 ( .INP(n7356), .ZN(n7231) );
  INVX0 U7320 ( .INP(n7356), .ZN(n7232) );
  INVX0 U7321 ( .INP(n7350), .ZN(n7233) );
  INVX0 U7322 ( .INP(n7351), .ZN(n7234) );
  INVX0 U7323 ( .INP(n7352), .ZN(n7235) );
  INVX0 U7324 ( .INP(n7349), .ZN(n7236) );
  INVX0 U7325 ( .INP(n7334), .ZN(n7237) );
  INVX0 U7326 ( .INP(n7347), .ZN(n7238) );
  INVX0 U7327 ( .INP(n7339), .ZN(n7239) );
  INVX0 U7328 ( .INP(n7339), .ZN(n7240) );
  INVX0 U7329 ( .INP(n7339), .ZN(n7241) );
  INVX0 U7330 ( .INP(n7339), .ZN(n7242) );
  INVX0 U7331 ( .INP(n7339), .ZN(n7243) );
  INVX0 U7332 ( .INP(n7339), .ZN(n7244) );
  INVX0 U7333 ( .INP(n7338), .ZN(n7245) );
  INVX0 U7334 ( .INP(n7338), .ZN(n7246) );
  INVX0 U7335 ( .INP(n7338), .ZN(n7247) );
  INVX0 U7336 ( .INP(n7338), .ZN(n7248) );
  INVX0 U7337 ( .INP(n7338), .ZN(n7249) );
  INVX0 U7338 ( .INP(n7338), .ZN(n7250) );
  INVX0 U7339 ( .INP(n7337), .ZN(n7251) );
  INVX0 U7340 ( .INP(n7337), .ZN(n7252) );
  INVX0 U7341 ( .INP(n7337), .ZN(n7253) );
  INVX0 U7342 ( .INP(n7337), .ZN(n7254) );
  INVX0 U7343 ( .INP(n7337), .ZN(n7255) );
  INVX0 U7344 ( .INP(n7337), .ZN(n7256) );
  INVX0 U7345 ( .INP(n7353), .ZN(n7257) );
  INVX0 U7346 ( .INP(n7343), .ZN(n7258) );
  INVX0 U7347 ( .INP(n7350), .ZN(n7259) );
  INVX0 U7348 ( .INP(n7346), .ZN(n7260) );
  INVX0 U7349 ( .INP(n7349), .ZN(n7261) );
  INVX0 U7350 ( .INP(n7357), .ZN(n7262) );
  INVX0 U7351 ( .INP(n7338), .ZN(n7263) );
  INVX0 U7352 ( .INP(n7342), .ZN(n7264) );
  INVX0 U7353 ( .INP(n7343), .ZN(n7265) );
  INVX0 U7354 ( .INP(n7341), .ZN(n7266) );
  INVX0 U7355 ( .INP(n7358), .ZN(n7267) );
  INVX0 U7356 ( .INP(n7354), .ZN(n7268) );
  INVX0 U7357 ( .INP(n7345), .ZN(n7269) );
  INVX0 U7358 ( .INP(n7340), .ZN(n7270) );
  INVX0 U7359 ( .INP(n7357), .ZN(n7271) );
  INVX0 U7360 ( .INP(n7356), .ZN(n7272) );
  INVX0 U7361 ( .INP(n7337), .ZN(n7273) );
  INVX0 U7362 ( .INP(n7344), .ZN(n7274) );
  INVX0 U7363 ( .INP(n7346), .ZN(n7275) );
  INVX0 U7364 ( .INP(n7334), .ZN(n7276) );
  INVX0 U7365 ( .INP(n7335), .ZN(n7277) );
  INVX0 U7366 ( .INP(n7336), .ZN(n7278) );
  INVX0 U7367 ( .INP(n7337), .ZN(n7279) );
  INVX0 U7368 ( .INP(n7348), .ZN(n7280) );
  INVX0 U7369 ( .INP(n7358), .ZN(n7281) );
  INVX0 U7370 ( .INP(n7341), .ZN(n7282) );
  INVX0 U7371 ( .INP(n7350), .ZN(n7283) );
  INVX0 U7372 ( .INP(n7334), .ZN(n7284) );
  INVX0 U7373 ( .INP(n7345), .ZN(n7285) );
  INVX0 U7374 ( .INP(n7357), .ZN(n7286) );
  INVX0 U7375 ( .INP(n7335), .ZN(n7287) );
  INVX0 U7376 ( .INP(n7340), .ZN(n7288) );
  INVX0 U7377 ( .INP(n7336), .ZN(n7289) );
  INVX0 U7378 ( .INP(n7347), .ZN(n7290) );
  INVX0 U7379 ( .INP(n7340), .ZN(n7291) );
  INVX0 U7380 ( .INP(n7344), .ZN(n7292) );
  INVX0 U7381 ( .INP(n7336), .ZN(n7293) );
  INVX0 U7382 ( .INP(n7336), .ZN(n7294) );
  INVX0 U7383 ( .INP(n7336), .ZN(n7295) );
  INVX0 U7384 ( .INP(n7336), .ZN(n7296) );
  INVX0 U7385 ( .INP(n7336), .ZN(n7297) );
  INVX0 U7386 ( .INP(n7336), .ZN(n7298) );
  INVX0 U7387 ( .INP(n7335), .ZN(n7299) );
  INVX0 U7388 ( .INP(n7335), .ZN(n7300) );
  INVX0 U7389 ( .INP(n7335), .ZN(n7301) );
  INVX0 U7390 ( .INP(n7335), .ZN(n7302) );
  INVX0 U7391 ( .INP(n7335), .ZN(n7303) );
  INVX0 U7392 ( .INP(n7335), .ZN(n7304) );
  INVX0 U7393 ( .INP(n7334), .ZN(n7305) );
  INVX0 U7394 ( .INP(n7334), .ZN(n7306) );
  INVX0 U7395 ( .INP(n7334), .ZN(n7307) );
  INVX0 U7396 ( .INP(n7334), .ZN(n7308) );
  INVX0 U7397 ( .INP(n7334), .ZN(n7309) );
  INVX0 U7398 ( .INP(n7334), .ZN(n7310) );
  INVX0 U7399 ( .INP(n7356), .ZN(n7311) );
  INVX0 U7400 ( .INP(n7339), .ZN(n7312) );
  INVX0 U7401 ( .INP(n7350), .ZN(n7313) );
  INVX0 U7402 ( .INP(n7346), .ZN(n7314) );
  INVX0 U7403 ( .INP(n7349), .ZN(n7315) );
  INVX0 U7404 ( .INP(n7341), .ZN(n7316) );
  INVX0 U7405 ( .INP(n7336), .ZN(n7317) );
  INVX0 U7406 ( .INP(n7342), .ZN(n7318) );
  INVX0 U7407 ( .INP(n7338), .ZN(n7319) );
  INVX0 U7408 ( .INP(n7339), .ZN(n7320) );
  INVX0 U7409 ( .INP(n7342), .ZN(n7321) );
  INVX0 U7410 ( .INP(n7343), .ZN(n7322) );
  INVX0 U7411 ( .INP(n7345), .ZN(n7323) );
  INVX0 U7412 ( .INP(n7346), .ZN(n7324) );
  INVX0 U7413 ( .INP(n7338), .ZN(n7325) );
  INVX0 U7414 ( .INP(n7358), .ZN(n7326) );
  INVX0 U7415 ( .INP(n7353), .ZN(n7327) );
  INVX0 U7416 ( .INP(n7340), .ZN(n7328) );
  INVX0 U7417 ( .INP(n7355), .ZN(n7329) );
  INVX0 U7418 ( .INP(n7340), .ZN(n7330) );
  INVX0 U7419 ( .INP(n7356), .ZN(n7331) );
  INVX0 U7420 ( .INP(n7355), .ZN(n7332) );
  INVX0 U7421 ( .INP(n7354), .ZN(n7333) );
  INVX0 U7422 ( .INP(rst), .ZN(n7358) );
endmodule


module RFSM_addrbits8_depth128 ( empty, rden, rdaddr, rdptr, sync_wrptr, 
        remove, clk_out, rst, sync_flush_BAR );
  output [7:0] rdaddr;
  output [8:0] rdptr;
  input [8:0] sync_wrptr;
  input remove, clk_out, rst, sync_flush_BAR;
  output empty, rden;
  wire   sync_flush, \rbin[8] , N12, N43, N44, N45, N46, N47, N48, N49, N50,
         N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, n12, n13, n14,
         \add_19/carry[8] , \add_19/carry[7] , \add_19/carry[6] ,
         \add_19/carry[5] , \add_19/carry[4] , \add_19/carry[3] ,
         \add_19/carry[2] , \add_19/carry[1] , n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27;
  wire   [8:0] rbinnext;
  wire   [7:0] rgraynext;
  wire   [1:0] next_state;
  wire   [1:0] current_state;
  assign sync_flush = sync_flush_BAR;

  DFFARX1 \rbin_reg[0]  ( .D(N44), .CLK(clk_out), .RSTB(n5), .Q(rdaddr[0]) );
  DFFASX1 empty_reg ( .D(N43), .CLK(clk_out), .SETB(n6), .Q(empty), .QN(n4) );
  DFFARX1 \current_state_reg[1]  ( .D(next_state[1]), .CLK(clk_out), .RSTB(n5), 
        .Q(current_state[1]) );
  DFFARX1 \current_state_reg[0]  ( .D(next_state[0]), .CLK(clk_out), .RSTB(n5), 
        .Q(current_state[0]) );
  DFFARX1 \rbin_reg[8]  ( .D(N52), .CLK(clk_out), .RSTB(n5), .Q(\rbin[8] ) );
  DFFARX1 \rbin_reg[1]  ( .D(N45), .CLK(clk_out), .RSTB(n5), .Q(rdaddr[1]) );
  DFFARX1 \rbin_reg[2]  ( .D(N46), .CLK(clk_out), .RSTB(n5), .Q(rdaddr[2]) );
  DFFARX1 \rbin_reg[3]  ( .D(N47), .CLK(clk_out), .RSTB(n5), .Q(rdaddr[3]) );
  DFFARX1 \rbin_reg[4]  ( .D(N48), .CLK(clk_out), .RSTB(n5), .Q(rdaddr[4]) );
  DFFARX1 \rbin_reg[5]  ( .D(N49), .CLK(clk_out), .RSTB(n5), .Q(rdaddr[5]) );
  DFFARX1 \rbin_reg[6]  ( .D(N50), .CLK(clk_out), .RSTB(n5), .Q(rdaddr[6]) );
  DFFARX1 \rbin_reg[7]  ( .D(N51), .CLK(clk_out), .RSTB(n5), .Q(rdaddr[7]) );
  DFFARX1 rden_reg ( .D(next_state[0]), .CLK(clk_out), .RSTB(n6), .Q(rden) );
  DFFARX1 \rdptr_reg[7]  ( .D(N60), .CLK(clk_out), .RSTB(n6), .Q(rdptr[7]) );
  DFFARX1 \rdptr_reg[6]  ( .D(N59), .CLK(clk_out), .RSTB(n6), .Q(rdptr[6]) );
  DFFARX1 \rdptr_reg[5]  ( .D(N58), .CLK(clk_out), .RSTB(n6), .Q(rdptr[5]) );
  DFFARX1 \rdptr_reg[4]  ( .D(N57), .CLK(clk_out), .RSTB(n6), .Q(rdptr[4]) );
  DFFARX1 \rdptr_reg[3]  ( .D(N56), .CLK(clk_out), .RSTB(n6), .Q(rdptr[3]) );
  DFFARX1 \rdptr_reg[2]  ( .D(N55), .CLK(clk_out), .RSTB(n6), .Q(rdptr[2]) );
  DFFARX1 \rdptr_reg[1]  ( .D(N54), .CLK(clk_out), .RSTB(n6), .Q(rdptr[1]) );
  DFFARX1 \rdptr_reg[0]  ( .D(N53), .CLK(clk_out), .RSTB(n5), .Q(rdptr[0]) );
  AO22X1 U12 ( .IN1(next_state[0]), .IN2(rgraynext[7]), .IN3(rdptr[7]), .IN4(
        next_state[1]), .Q(N60) );
  XOR2X1 U13 ( .IN1(rbinnext[7]), .IN2(rbinnext[8]), .Q(rgraynext[7]) );
  AO22X1 U14 ( .IN1(next_state[0]), .IN2(rgraynext[6]), .IN3(rdptr[6]), .IN4(
        next_state[1]), .Q(N59) );
  XOR2X1 U15 ( .IN1(rbinnext[6]), .IN2(rbinnext[7]), .Q(rgraynext[6]) );
  AO22X1 U16 ( .IN1(next_state[0]), .IN2(rgraynext[5]), .IN3(rdptr[5]), .IN4(
        next_state[1]), .Q(N58) );
  XOR2X1 U17 ( .IN1(rbinnext[5]), .IN2(rbinnext[6]), .Q(rgraynext[5]) );
  AO22X1 U18 ( .IN1(next_state[0]), .IN2(rgraynext[4]), .IN3(rdptr[4]), .IN4(
        next_state[1]), .Q(N57) );
  XOR2X1 U19 ( .IN1(rbinnext[4]), .IN2(rbinnext[5]), .Q(rgraynext[4]) );
  AO22X1 U20 ( .IN1(next_state[0]), .IN2(rgraynext[3]), .IN3(rdptr[3]), .IN4(
        next_state[1]), .Q(N56) );
  XOR2X1 U21 ( .IN1(rbinnext[3]), .IN2(rbinnext[4]), .Q(rgraynext[3]) );
  AO22X1 U22 ( .IN1(next_state[0]), .IN2(rgraynext[2]), .IN3(rdptr[2]), .IN4(
        next_state[1]), .Q(N55) );
  XOR2X1 U23 ( .IN1(rbinnext[2]), .IN2(rbinnext[3]), .Q(rgraynext[2]) );
  AO22X1 U24 ( .IN1(next_state[0]), .IN2(rgraynext[1]), .IN3(rdptr[1]), .IN4(
        next_state[1]), .Q(N54) );
  XOR2X1 U25 ( .IN1(rbinnext[1]), .IN2(rbinnext[2]), .Q(rgraynext[1]) );
  AO22X1 U26 ( .IN1(next_state[0]), .IN2(rgraynext[0]), .IN3(rdptr[0]), .IN4(
        next_state[1]), .Q(N53) );
  XOR2X1 U27 ( .IN1(rbinnext[0]), .IN2(rbinnext[1]), .Q(rgraynext[0]) );
  AO22X1 U28 ( .IN1(next_state[0]), .IN2(rbinnext[8]), .IN3(\rbin[8] ), .IN4(
        next_state[1]), .Q(N52) );
  AO22X1 U29 ( .IN1(next_state[0]), .IN2(rbinnext[7]), .IN3(rdaddr[7]), .IN4(
        next_state[1]), .Q(N51) );
  AO22X1 U30 ( .IN1(next_state[0]), .IN2(rbinnext[6]), .IN3(rdaddr[6]), .IN4(
        next_state[1]), .Q(N50) );
  AO22X1 U31 ( .IN1(next_state[0]), .IN2(rbinnext[5]), .IN3(rdaddr[5]), .IN4(
        next_state[1]), .Q(N49) );
  AO22X1 U32 ( .IN1(next_state[0]), .IN2(rbinnext[4]), .IN3(rdaddr[4]), .IN4(
        next_state[1]), .Q(N48) );
  AO22X1 U33 ( .IN1(next_state[0]), .IN2(rbinnext[3]), .IN3(rdaddr[3]), .IN4(
        next_state[1]), .Q(N47) );
  AO22X1 U34 ( .IN1(next_state[0]), .IN2(rbinnext[2]), .IN3(rdaddr[2]), .IN4(
        next_state[1]), .Q(N46) );
  AO22X1 U35 ( .IN1(next_state[0]), .IN2(rbinnext[1]), .IN3(rdaddr[1]), .IN4(
        next_state[1]), .Q(N45) );
  AO22X1 U36 ( .IN1(next_state[0]), .IN2(rbinnext[0]), .IN3(rdaddr[0]), .IN4(
        next_state[1]), .Q(N44) );
  OAI22X1 U39 ( .IN1(N12), .IN2(current_state[0]), .IN3(n13), .IN4(
        current_state[1]), .QN(n12) );
  AND2X1 U40 ( .IN1(current_state[0]), .IN2(N12), .Q(n13) );
  AND3X1 U41 ( .IN1(n14), .IN2(sync_flush), .IN3(N12), .Q(next_state[0]) );
  XOR2X1 U42 ( .IN1(current_state[1]), .IN2(current_state[0]), .Q(n14) );
  AO21X1 U3 ( .IN1(n23), .IN2(rgraynext[1]), .IN3(n11), .Q(n18) );
  INVX0 U4 ( .INP(rgraynext[0]), .ZN(n24) );
  INVX0 U5 ( .INP(rgraynext[1]), .ZN(n25) );
  NAND3X0 U6 ( .IN1(n1), .IN2(n2), .IN3(n3), .QN(N43) );
  NOR2X0 U7 ( .IN1(n27), .IN2(rdaddr[7]), .QN(n1) );
  OR4X1 U8 ( .IN1(n22), .IN2(n21), .IN3(n20), .IN4(n19), .Q(n2) );
  OR2X1 U9 ( .IN1(next_state[1]), .IN2(next_state[0]), .Q(n3) );
  AND2X1 U10 ( .IN1(remove), .IN2(n4), .Q(N12) );
  AND2X1 U11 ( .IN1(n12), .IN2(sync_flush), .Q(next_state[1]) );
  NBUFFX2 U37 ( .INP(rst), .Z(n5) );
  NBUFFX2 U38 ( .INP(rst), .Z(n6) );
  INVX0 U43 ( .INP(sync_wrptr[1]), .ZN(n23) );
  XOR2X1 U44 ( .IN1(\rbin[8] ), .IN2(\add_19/carry[8] ), .Q(rbinnext[8]) );
  AND2X1 U45 ( .IN1(rdaddr[7]), .IN2(\add_19/carry[7] ), .Q(\add_19/carry[8] )
         );
  XOR2X1 U46 ( .IN1(rdaddr[7]), .IN2(\add_19/carry[7] ), .Q(rbinnext[7]) );
  AND2X1 U47 ( .IN1(rdaddr[6]), .IN2(\add_19/carry[6] ), .Q(\add_19/carry[7] )
         );
  XOR2X1 U48 ( .IN1(rdaddr[6]), .IN2(\add_19/carry[6] ), .Q(rbinnext[6]) );
  AND2X1 U49 ( .IN1(rdaddr[5]), .IN2(\add_19/carry[5] ), .Q(\add_19/carry[6] )
         );
  XOR2X1 U50 ( .IN1(rdaddr[5]), .IN2(\add_19/carry[5] ), .Q(rbinnext[5]) );
  AND2X1 U51 ( .IN1(rdaddr[4]), .IN2(\add_19/carry[4] ), .Q(\add_19/carry[5] )
         );
  XOR2X1 U52 ( .IN1(rdaddr[4]), .IN2(\add_19/carry[4] ), .Q(rbinnext[4]) );
  AND2X1 U53 ( .IN1(rdaddr[3]), .IN2(\add_19/carry[3] ), .Q(\add_19/carry[4] )
         );
  XOR2X1 U54 ( .IN1(rdaddr[3]), .IN2(\add_19/carry[3] ), .Q(rbinnext[3]) );
  AND2X1 U55 ( .IN1(rdaddr[2]), .IN2(\add_19/carry[2] ), .Q(\add_19/carry[3] )
         );
  XOR2X1 U56 ( .IN1(rdaddr[2]), .IN2(\add_19/carry[2] ), .Q(rbinnext[2]) );
  AND2X1 U57 ( .IN1(rdaddr[1]), .IN2(\add_19/carry[1] ), .Q(\add_19/carry[2] )
         );
  XOR2X1 U58 ( .IN1(rdaddr[1]), .IN2(\add_19/carry[1] ), .Q(rbinnext[1]) );
  AND2X1 U59 ( .IN1(rdaddr[0]), .IN2(N12), .Q(\add_19/carry[1] ) );
  XOR2X1 U60 ( .IN1(rdaddr[0]), .IN2(N12), .Q(rbinnext[0]) );
  XNOR2X1 U61 ( .IN1(sync_wrptr[8]), .IN2(rbinnext[8]), .Q(n10) );
  XNOR2X1 U62 ( .IN1(sync_wrptr[7]), .IN2(rgraynext[7]), .Q(n9) );
  XNOR2X1 U63 ( .IN1(sync_wrptr[6]), .IN2(rgraynext[6]), .Q(n8) );
  XNOR2X1 U64 ( .IN1(sync_wrptr[5]), .IN2(rgraynext[5]), .Q(n7) );
  NAND4X0 U65 ( .IN1(n10), .IN2(n9), .IN3(n8), .IN4(n7), .QN(n22) );
  NOR2X0 U66 ( .IN1(n24), .IN2(sync_wrptr[0]), .QN(n11) );
  AND2X1 U67 ( .IN1(sync_wrptr[0]), .IN2(n24), .Q(n15) );
  OA22X1 U68 ( .IN1(sync_wrptr[1]), .IN2(n15), .IN3(n15), .IN4(n25), .Q(n17)
         );
  XOR2X1 U69 ( .IN1(sync_wrptr[2]), .IN2(rgraynext[2]), .Q(n16) );
  OR3X1 U70 ( .IN1(n18), .IN2(n17), .IN3(n16), .Q(n21) );
  XOR2X1 U71 ( .IN1(sync_wrptr[3]), .IN2(rgraynext[3]), .Q(n20) );
  XOR2X1 U72 ( .IN1(sync_wrptr[4]), .IN2(rgraynext[4]), .Q(n19) );
  AND4X1 U73 ( .IN1(rdaddr[6]), .IN2(rdaddr[5]), .IN3(rdaddr[4]), .IN4(
        rdaddr[0]), .Q(n26) );
  AND4X1 U74 ( .IN1(rdaddr[3]), .IN2(rdaddr[2]), .IN3(rdaddr[1]), .IN4(n26), 
        .Q(n27) );
endmodule


module WFSM_addrbits8_depth128 ( full, wraddr, wrptr, sync_rdptr, insert, 
        flush, clk_in, rst, wren_BAR );
  output [7:0] wraddr;
  output [8:0] wrptr;
  input [8:0] sync_rdptr;
  input insert, flush, clk_in, rst;
  output full, wren_BAR;
  wire   \wbin[8] , N10, N12, N13, \next_state[1] , N42, N43, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, \add_19/carry[8] ,
         \add_19/carry[7] , \add_19/carry[6] , \add_19/carry[5] ,
         \add_19/carry[4] , \add_19/carry[3] , \add_19/carry[2] ,
         \add_19/carry[1] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n37, n38, n39, n40, n41, n42, n43, n45, n46;
  wire   [8:0] wbinnext;
  wire   [7:0] wgraynext;
  wire   [1:0] current_state;

  DFFARX1 \wbin_reg[0]  ( .D(n36), .CLK(clk_in), .RSTB(n3), .Q(wraddr[0]) );
  DFFARX1 full_reg ( .D(N43), .CLK(clk_in), .RSTB(n3), .Q(full), .QN(n1) );
  DFFARX1 \current_state_reg[1]  ( .D(\next_state[1] ), .CLK(clk_in), .RSTB(n3), .Q(current_state[1]) );
  DFFARX1 \current_state_reg[0]  ( .D(n46), .CLK(clk_in), .RSTB(n3), .Q(
        current_state[0]) );
  DFFARX1 wren_reg ( .D(N42), .CLK(clk_in), .RSTB(n3), .QN(wren_BAR) );
  DFFARX1 \wbin_reg[7]  ( .D(n28), .CLK(clk_in), .RSTB(n3), .Q(wraddr[7]) );
  DFFARX1 \wbin_reg[1]  ( .D(n34), .CLK(clk_in), .RSTB(n3), .Q(wraddr[1]) );
  DFFARX1 \wbin_reg[2]  ( .D(n33), .CLK(clk_in), .RSTB(n3), .Q(wraddr[2]) );
  DFFARX1 \wbin_reg[3]  ( .D(n32), .CLK(clk_in), .RSTB(n3), .Q(wraddr[3]) );
  DFFARX1 \wbin_reg[4]  ( .D(n31), .CLK(clk_in), .RSTB(n3), .Q(wraddr[4]) );
  DFFARX1 \wbin_reg[5]  ( .D(n30), .CLK(clk_in), .RSTB(n2), .Q(wraddr[5]) );
  DFFARX1 \wbin_reg[6]  ( .D(n29), .CLK(clk_in), .RSTB(n2), .Q(wraddr[6]) );
  DFFARX1 \wbin_reg[8]  ( .D(n35), .CLK(clk_in), .RSTB(n2), .Q(\wbin[8] ) );
  DFFARX1 \wrptr_reg[0]  ( .D(n27), .CLK(clk_in), .RSTB(n2), .Q(wrptr[0]) );
  DFFARX1 \wrptr_reg[1]  ( .D(n26), .CLK(clk_in), .RSTB(n2), .Q(wrptr[1]) );
  DFFARX1 \wrptr_reg[2]  ( .D(n25), .CLK(clk_in), .RSTB(n2), .Q(wrptr[2]) );
  DFFARX1 \wrptr_reg[3]  ( .D(n24), .CLK(clk_in), .RSTB(n2), .Q(wrptr[3]) );
  DFFARX1 \wrptr_reg[4]  ( .D(n23), .CLK(clk_in), .RSTB(n2), .Q(wrptr[4]) );
  DFFARX1 \wrptr_reg[5]  ( .D(n22), .CLK(clk_in), .RSTB(n2), .Q(wrptr[5]) );
  DFFARX1 \wrptr_reg[6]  ( .D(n21), .CLK(clk_in), .RSTB(n2), .Q(wrptr[6]) );
  DFFARX1 \wrptr_reg[7]  ( .D(n20), .CLK(clk_in), .RSTB(n2), .Q(wrptr[7]) );
  DFFARX1 \wrptr_reg[8]  ( .D(n19), .CLK(clk_in), .RSTB(n2), .Q(wrptr[8]) );
  AO22X1 U15 ( .IN1(wrptr[8]), .IN2(n13), .IN3(N42), .IN4(wbinnext[8]), .Q(n19) );
  AO22X1 U16 ( .IN1(wrptr[7]), .IN2(n13), .IN3(N42), .IN4(n14), .Q(n20) );
  AO22X1 U17 ( .IN1(wrptr[6]), .IN2(n13), .IN3(N42), .IN4(wgraynext[6]), .Q(
        n21) );
  XOR2X1 U18 ( .IN1(wbinnext[6]), .IN2(wbinnext[7]), .Q(wgraynext[6]) );
  AO22X1 U19 ( .IN1(wrptr[5]), .IN2(n13), .IN3(N42), .IN4(wgraynext[5]), .Q(
        n22) );
  XOR2X1 U20 ( .IN1(wbinnext[5]), .IN2(wbinnext[6]), .Q(wgraynext[5]) );
  AO22X1 U21 ( .IN1(wrptr[4]), .IN2(n13), .IN3(N42), .IN4(wgraynext[4]), .Q(
        n23) );
  XOR2X1 U22 ( .IN1(wbinnext[4]), .IN2(wbinnext[5]), .Q(wgraynext[4]) );
  AO22X1 U23 ( .IN1(wrptr[3]), .IN2(n13), .IN3(N42), .IN4(wgraynext[3]), .Q(
        n24) );
  XOR2X1 U24 ( .IN1(wbinnext[3]), .IN2(wbinnext[4]), .Q(wgraynext[3]) );
  AO22X1 U25 ( .IN1(wrptr[2]), .IN2(n13), .IN3(N42), .IN4(wgraynext[2]), .Q(
        n25) );
  XOR2X1 U26 ( .IN1(wbinnext[2]), .IN2(wbinnext[3]), .Q(wgraynext[2]) );
  AO22X1 U27 ( .IN1(wrptr[1]), .IN2(n13), .IN3(N42), .IN4(wgraynext[1]), .Q(
        n26) );
  XOR2X1 U28 ( .IN1(wbinnext[1]), .IN2(wbinnext[2]), .Q(wgraynext[1]) );
  AO22X1 U29 ( .IN1(wrptr[0]), .IN2(n13), .IN3(N42), .IN4(wgraynext[0]), .Q(
        n27) );
  XOR2X1 U30 ( .IN1(wbinnext[0]), .IN2(wbinnext[1]), .Q(wgraynext[0]) );
  AO22X1 U31 ( .IN1(wraddr[7]), .IN2(n13), .IN3(N42), .IN4(wbinnext[7]), .Q(
        n28) );
  AO22X1 U32 ( .IN1(wraddr[6]), .IN2(n13), .IN3(N42), .IN4(wbinnext[6]), .Q(
        n29) );
  AO22X1 U33 ( .IN1(wraddr[5]), .IN2(n13), .IN3(N42), .IN4(wbinnext[5]), .Q(
        n30) );
  AO22X1 U34 ( .IN1(wraddr[4]), .IN2(n13), .IN3(N42), .IN4(wbinnext[4]), .Q(
        n31) );
  AO22X1 U35 ( .IN1(wraddr[3]), .IN2(n13), .IN3(N42), .IN4(wbinnext[3]), .Q(
        n32) );
  AO22X1 U36 ( .IN1(wraddr[2]), .IN2(n13), .IN3(N42), .IN4(wbinnext[2]), .Q(
        n33) );
  AO22X1 U37 ( .IN1(wraddr[1]), .IN2(n13), .IN3(N42), .IN4(wbinnext[1]), .Q(
        n34) );
  AO22X1 U38 ( .IN1(\wbin[8] ), .IN2(n13), .IN3(N42), .IN4(wbinnext[8]), .Q(
        n35) );
  AO22X1 U39 ( .IN1(wraddr[0]), .IN2(n13), .IN3(N42), .IN4(wbinnext[0]), .Q(
        n36) );
  AND3X1 U41 ( .IN1(n45), .IN2(n4), .IN3(n17), .Q(\next_state[1] ) );
  AO21X1 U42 ( .IN1(N12), .IN2(n18), .IN3(N13), .Q(n15) );
  XOR2X1 U43 ( .IN1(sync_rdptr[7]), .IN2(n14), .Q(n18) );
  XOR2X1 U44 ( .IN1(wbinnext[7]), .IN2(wbinnext[8]), .Q(n14) );
  NAND3X0 U45 ( .IN1(n17), .IN2(n4), .IN3(N10), .QN(n16) );
  AO21X1 U3 ( .IN1(n39), .IN2(wgraynext[1]), .IN3(n5), .Q(n8) );
  INVX0 U4 ( .INP(wgraynext[0]), .ZN(n40) );
  INVX0 U5 ( .INP(wgraynext[1]), .ZN(n41) );
  INVX0 U6 ( .INP(n16), .ZN(n46) );
  NOR2X0 U7 ( .IN1(n16), .IN2(n15), .QN(N42) );
  AO21X1 U8 ( .IN1(n46), .IN2(n15), .IN3(\next_state[1] ), .Q(n13) );
  OA21X1 U9 ( .IN1(\next_state[1] ), .IN2(n46), .IN3(n15), .Q(N43) );
  INVX0 U10 ( .INP(N10), .ZN(n45) );
  AND2X1 U11 ( .IN1(insert), .IN2(n1), .Q(N10) );
  AND2X1 U12 ( .IN1(wraddr[1]), .IN2(\add_19/carry[1] ), .Q(\add_19/carry[2] )
         );
  AND2X1 U13 ( .IN1(wraddr[3]), .IN2(\add_19/carry[3] ), .Q(\add_19/carry[4] )
         );
  XOR2X1 U14 ( .IN1(wraddr[1]), .IN2(\add_19/carry[1] ), .Q(wbinnext[1]) );
  XOR2X1 U40 ( .IN1(wraddr[3]), .IN2(\add_19/carry[3] ), .Q(wbinnext[3]) );
  AND4X1 U46 ( .IN1(wraddr[3]), .IN2(wraddr[2]), .IN3(wraddr[1]), .IN4(n42), 
        .Q(n43) );
  NAND2X1 U47 ( .IN1(current_state[1]), .IN2(current_state[0]), .QN(n17) );
  NBUFFX2 U48 ( .INP(rst), .Z(n2) );
  NBUFFX2 U49 ( .INP(rst), .Z(n3) );
  INVX0 U50 ( .INP(sync_rdptr[1]), .ZN(n39) );
  INVX0 U51 ( .INP(flush), .ZN(n4) );
  XOR2X1 U52 ( .IN1(\wbin[8] ), .IN2(\add_19/carry[8] ), .Q(wbinnext[8]) );
  AND2X1 U53 ( .IN1(wraddr[7]), .IN2(\add_19/carry[7] ), .Q(\add_19/carry[8] )
         );
  XOR2X1 U54 ( .IN1(wraddr[7]), .IN2(\add_19/carry[7] ), .Q(wbinnext[7]) );
  AND2X1 U55 ( .IN1(wraddr[6]), .IN2(\add_19/carry[6] ), .Q(\add_19/carry[7] )
         );
  XOR2X1 U56 ( .IN1(wraddr[6]), .IN2(\add_19/carry[6] ), .Q(wbinnext[6]) );
  AND2X1 U57 ( .IN1(wraddr[5]), .IN2(\add_19/carry[5] ), .Q(\add_19/carry[6] )
         );
  XOR2X1 U58 ( .IN1(wraddr[5]), .IN2(\add_19/carry[5] ), .Q(wbinnext[5]) );
  AND2X1 U59 ( .IN1(wraddr[4]), .IN2(\add_19/carry[4] ), .Q(\add_19/carry[5] )
         );
  XOR2X1 U60 ( .IN1(wraddr[4]), .IN2(\add_19/carry[4] ), .Q(wbinnext[4]) );
  AND2X1 U61 ( .IN1(wraddr[2]), .IN2(\add_19/carry[2] ), .Q(\add_19/carry[3] )
         );
  XOR2X1 U62 ( .IN1(wraddr[2]), .IN2(\add_19/carry[2] ), .Q(wbinnext[2]) );
  AND2X1 U63 ( .IN1(wraddr[0]), .IN2(N10), .Q(\add_19/carry[1] ) );
  XOR2X1 U64 ( .IN1(wraddr[0]), .IN2(N10), .Q(wbinnext[0]) );
  XOR2X1 U65 ( .IN1(sync_rdptr[2]), .IN2(wgraynext[2]), .Q(n10) );
  XOR2X1 U66 ( .IN1(sync_rdptr[3]), .IN2(wgraynext[3]), .Q(n9) );
  NOR2X0 U67 ( .IN1(n40), .IN2(sync_rdptr[0]), .QN(n5) );
  AND2X1 U68 ( .IN1(sync_rdptr[0]), .IN2(n40), .Q(n6) );
  OA22X1 U69 ( .IN1(sync_rdptr[1]), .IN2(n6), .IN3(n6), .IN4(n41), .Q(n7) );
  OR4X1 U70 ( .IN1(n10), .IN2(n9), .IN3(n8), .IN4(n7), .Q(n38) );
  XOR2X1 U71 ( .IN1(sync_rdptr[6]), .IN2(wgraynext[6]), .Q(n37) );
  XOR2X1 U72 ( .IN1(sync_rdptr[4]), .IN2(wgraynext[4]), .Q(n12) );
  XOR2X1 U73 ( .IN1(sync_rdptr[5]), .IN2(wgraynext[5]), .Q(n11) );
  NOR4X0 U74 ( .IN1(n38), .IN2(n37), .IN3(n12), .IN4(n11), .QN(N12) );
  AND4X1 U75 ( .IN1(wraddr[6]), .IN2(wraddr[5]), .IN3(wraddr[4]), .IN4(
        wraddr[0]), .Q(n42) );
  OR2X1 U76 ( .IN1(n43), .IN2(wraddr[7]), .Q(N13) );
endmodule


module fifo ( dataOut, full, empty, dataIn, insert, flush, clk_in, rst, remove, 
        clk_out );
  output [31:0] dataOut;
  input [31:0] dataIn;
  input insert, flush, clk_in, rst, remove, clk_out;
  output full, empty;
  wire   sync_flush, wren, rden;
  wire   [8:0] sync_rdptr;
  wire   [8:0] rdptr;
  wire   [8:0] sync_wrptr;
  wire   [8:0] wrptr;
  wire   [7:0] wraddr;
  wire   [7:0] rdaddr;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;

  read_sync_addrbits8 r2w_uut ( .clk_out(clk_out), .rst(rst), .rdptr({1'b0, 
        rdptr[7:0]}), .sync_rdptr({SYNOPSYS_UNCONNECTED__0, sync_rdptr[7:0]}), 
        .sync_flush_BAR(sync_flush) );
  write_sync_addrbits8 w2r_uut ( .clk_in(clk_in), .rst(rst), .flush(flush), 
        .wrptr(wrptr), .sync_wrptr(sync_wrptr) );
  flush_sync flush_uut ( .clk_in(clk_in), .rst(rst), .flush(flush), 
        .sync_flush_BAR(sync_flush) );
  memory_datasize32_addrbits8_depth128 mem_uut ( .clk_in(clk_in), .flush(flush), .rst(rst), .clk_out(clk_out), .rden(rden), .rdaddr(rdaddr), .wraddr(wraddr), 
        .dataIn(dataIn), .dataOut(dataOut), .sync_flush_BAR(sync_flush), 
        .wren_BAR(wren) );
  RFSM_addrbits8_depth128 read_uut ( .empty(empty), .rden(rden), .rdaddr(
        rdaddr), .rdptr({SYNOPSYS_UNCONNECTED__1, rdptr[7:0]}), .sync_wrptr(
        sync_wrptr), .remove(remove), .clk_out(clk_out), .rst(rst), 
        .sync_flush_BAR(sync_flush) );
  WFSM_addrbits8_depth128 write_uut ( .full(full), .wraddr(wraddr), .wrptr(
        wrptr), .sync_rdptr({1'b0, sync_rdptr[7:0]}), .insert(insert), .flush(
        flush), .clk_in(clk_in), .rst(rst), .wren_BAR(wren) );
endmodule

